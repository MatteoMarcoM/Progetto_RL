//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "it"
//: property prefix = "_GG"
//: property title = "flipflopd.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
supply0 w6;    //: /sn:0 {0}(840,393)(840,354)(774,354){1}
reg [7:0] b;    //: /sn:0 {0}(#:254,-645)(254,-694){1}
//: {2}(#:256,-696)(352,-696)(352,-721){3}
//: {4}(254,-698)(#:254,-714){5}
//: {6}(#:252,-696)(137,-696)(137,-734){7}
supply0 w19;    //: /sn:0 {0}(177,3)(177,-16)(269,-16){1}
//: {2}(273,-16)(321,-16){3}
//: {4}(271,-18)(271,-26)(321,-26){5}
supply0 w21;    //: /sn:0 {0}(788,-353)(714,-353)(714,-345){1}
//: {2}(716,-343)(788,-343){3}
//: {4}(712,-343)(664,-343)(664,-326){5}
supply1 w1;    //: /sn:0 {0}(1104,-179)(1104,-169)(1062,-169)(1062,-223)(1095,-223){1}
reg clk;    //: /sn:0 {0}(1104,6)(1136,6)(1136,-54)(792,-54)(792,-226){1}
//: {2}(794,-228)(917,-228){3}
//: {4}(790,-228)(584,-228){5}
//: {6}(582,-230)(582,-385)(581,-385)(581,-584){7}
//: {8}(583,-586)(665,-586){9}
//: {10}(669,-586)(719,-586){11}
//: {12}(667,-584)(667,-530)(877,-530)(877,-582)(985,-582){13}
//: {14}(581,-588)(581,-663)(195,-663){15}
//: {16}(191,-663)(140,-663)(140,-419){17}
//: {18}(142,-417)(189,-417)(189,-372){19}
//: {20}(138,-417)(46,-417)(46,498)(767,498){21}
//: {22}(771,498)(819,498){23}
//: {24}(769,500)(769,613)(1304,613)(1304,497)(1353,497){25}
//: {26}(193,-661)(193,-645){27}
//: {28}(579,-586)(518,-586){29}
//: {30}(580,-228)(465,-228)(465,-76)(343,-76)(343,22){31}
reg [7:0] a;    //: /sn:0 {0}(#:683,-707)(683,-693){1}
//: {2}(#:685,-691)(768,-691)(768,-728){3}
//: {4}(#:681,-691)(574,-691)(574,-725){5}
//: {6}(683,-689)(683,-647)(#:719,-647){7}
reg [7:0] c;    //: /sn:0 {0}(#:962,-692)(962,-684){1}
//: {2}(#:964,-682)(1041,-682){3}
//: {4}(#:1045,-682)(1124,-682)(1124,-711){5}
//: {6}(1043,-684)(1043,-710){7}
//: {8}(962,-680)(962,-643)(#:985,-643){9}
wire [17:0] w16;    //: /sn:0 {0}(#:979,28)(816,28)(816,223){1}
//: {2}(818,225)(965,225){3}
//: {4}(969,225)(1117,225)(1117,189){5}
//: {6}(967,223)(#:967,148){7}
//: {8}(814,225)(725,225)(#:725,294){9}
wire [17:0] delta;    //: /sn:0 {0}(#:1478,475)(1552,475){1}
//: {2}(1556,475)(1691,475)(1691,415){3}
//: {4}(1554,473)(1554,424){5}
wire w4;    //: /sn:0 {0}(1058,480)(1058,501){1}
//: {2}(1060,503)(1103,503){3}
//: {4}(1058,505)(1058,567)(1796,567)(1796,427){5}
wire [7:0] w15;    //: /sn:0 {0}(#:839,-565)(839,-643)(#:809,-643){1}
wire w3;    //: /sn:0 {0}(568,320)(568,357)(608,357){1}
wire [17:0] w0;    //: /sn:0 {0}(#:1103,476)(1058,476){1}
//: {2}(1057,476)(991,476){3}
//: {4}(989,474)(989,425){5}
//: {6}(987,476)(#:944,476){7}
//: {8}(989,478)(989,520){9}
wire [7:0] w20;    //: /sn:0 {0}(#:250,-372)(#:250,-555){1}
wire [15:0] w23;    //: /sn:0 {0}(#:788,-363)(699,-363)(699,-390){1}
//: {2}(701,-392)(848,-392){3}
//: {4}(852,-392)(1052,-392)(1052,-460){5}
//: {6}(850,-394)(#:850,-425){7}
//: {8}(#:697,-392)(647,-392)(647,-427){9}
wire [7:0] w25;    //: /sn:0 {0}(#:246,-282)(246,-249){1}
//: {2}(248,-247)(380,-247)(380,-150)(#:339,-150){3}
//: {4}(246,-245)(#:246,-220){5}
wire [17:0] w8;    //: /sn:0 {0}(#:365,147)(365,210)(489,210){1}
//: {2}(493,210)(627,210){3}
//: {4}(631,210)(632,210)(#:632,294){5}
//: {6}(629,208)(629,135){7}
//: {8}(491,208)(491,142){9}
wire [17:0] w18;    //: /sn:0 {0}(#:917,-251)(899,-251)(899,-353)(#:794,-353){1}
wire [7:0] w17;    //: /sn:0 {0}(#:932,-495)(947,-495)(947,-533)(1085,-533)(1085,-639)(#:1075,-639){1}
wire [17:0] w22;    //: /sn:0 {0}(#:1095,-250)(1070,-250){1}
//: {2}(1068,-252)(1068,-289){3}
//: {4}(1068,-293)(1068,-334){5}
//: {6}(#:1066,-291)(981,-291)(981,-305){7}
//: {8}(1066,-250)(#:1042,-250){9}
wire [17:0] w11;    //: /sn:0 {0}(819,475)(677,475)(#:677,438){1}
wire [17:0] w12;    //: /sn:0 {0}(#:1104,29)(1269,29)(1269,-252)(#:1235,-252){1}
wire [17:0] w27;    //: /sn:0 {0}(#:366,22)(366,-26)(#:327,-26){1}
wire [17:0] w13;    //: /sn:0 {0}(#:1353,474)(#:1243,474){1}
wire w5;    //: /sn:0 {0}(1158,-287)(1158,-310)(1226,-310)(1226,-369){1}
wire w9;    //: /sn:0 {0}(1213,404)(1213,424)(1166,424)(1166,439){1}
wire [15:0] w26;    //: /sn:0 {0}(321,-36)(257,-36)(#:257,-80){1}
//: enddecls

  //: GROUND g4 (w6) @(840,399) /sn:0 /w:[ 0 ]
  //: joint g8 (w16) @(816, 225) /w:[ 2 1 8 -1 ]
  //: joint g61 (w23) @(699, -392) /w:[ 2 -1 8 1 ]
  //: LED g34 (w23) @(1052,-467) /sn:0 /w:[ 5 ] /type:3
  MyCOMPLEMENT2 g13 (.minus(w1), .In(w22), .Cout(w5), .Out(w12));   //: @(1096, -286) /sz:(138, 79) /sn:0 /p:[ Li0>1 Li1>0 To0<0 Ro0<1 ]
  //: LED g3 (w8) @(491,135) /sn:0 /w:[ 9 ] /type:3
  MYREGISTER8 g37 (.in(b), .Clk(clk), .out(w20));   //: @(177, -644) /sz:(106, 88) /R:3 /sn:0 /p:[ Ti0>0 Ti1>27 Bo0<1 ]
  //: LED g51 (w22) @(1068,-341) /sn:0 /w:[ 5 ] /type:3
  //: LED g55 (w0) @(989,527) /sn:0 /R:2 /w:[ 9 ] /type:1
  //: LED g58 (w8) @(629,128) /sn:0 /w:[ 7 ] /type:1
  //: joint g2 (w8) @(491, 210) /w:[ 2 8 1 -1 ]
  assign w4 = w0[17]; //: TAP g65 @(1058,474) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  //: joint g59 (w8) @(629, 210) /w:[ 4 6 3 -1 ]
  //: LED g1 (w16) @(967,141) /sn:0 /w:[ 7 ] /type:3
  //: LED g64 (w4) @(1796,420) /sn:0 /w:[ 5 ] /type:0
  MyCOMPLEMENT2 g11 (.minus(w4), .In(w0), .Cout(w9), .Out(w13));   //: @(1104, 440) /sz:(138, 79) /sn:0 /p:[ Li0>3 Li1>0 To0<1 Ro0<1 ]
  MYREGISTER18 g16 (.Clk(clk), .in(w13), .out(delta));   //: @(1354, 463) /sz:(123, 41) /sn:0 /p:[ Li0>25 Li1>0 Ro0<0 ]
  //: DIP g28 (c) @(962,-702) /sn:0 /w:[ 0 ] /st:5 /dn:1
  //: LED g10 (delta) @(1691,408) /sn:0 /w:[ 3 ] /type:1
  //: joint g50 (clk) @(582, -228) /w:[ 5 6 30 -1 ]
  //: LED g32 (c) @(1043,-717) /sn:0 /w:[ 7 ] /type:3
  //: DIP g27 (a) @(683,-717) /sn:0 /w:[ 0 ] /st:3 /dn:1
  //: joint g19 (clk) @(769, 498) /w:[ 22 -1 21 24 ]
  //: LED g69 (a) @(574,-732) /sn:0 /w:[ 5 ] /type:1
  MYREGISTER18 g6 (.in(w11), .Clk(clk), .out(w0));   //: @(820, 464) /sz:(123, 41) /sn:0 /p:[ Li0>0 Li1>23 Ro0<7 ]
  //: joint g38 (clk) @(581, -586) /w:[ 8 14 28 7 ]
  //: SWITCH g7 (clk) @(501,-586) /sn:0 /w:[ 29 ] /st:1 /dn:1
  //: joint g9 (clk) @(140, -417) /w:[ 18 17 20 -1 ]
  //: LED g53 (w5) @(1226,-376) /sn:0 /w:[ 1 ] /type:0
  //: joint g57 (w16) @(967, 225) /w:[ 4 6 3 -1 ]
  //: joint g71 (c) @(1043, -682) /w:[ 4 6 3 -1 ]
  //: joint g31 (a) @(683, -691) /w:[ 2 1 4 6 ]
  //: joint g15 (clk) @(792, -228) /w:[ 2 -1 4 1 ]
  //: VDD g20 (w1) @(1115,-179) /sn:0 /w:[ 0 ]
  //: LED g68 (b) @(137,-741) /sn:0 /w:[ 7 ] /type:1
  //: joint g67 (b) @(254, -696) /w:[ 2 4 6 1 ]
  //: joint g39 (w23) @(850, -392) /w:[ 4 6 3 -1 ]
  //: joint g43 (clk) @(193, -663) /w:[ 15 -1 16 26 ]
  //: joint g48 (w19) @(271, -16) /w:[ 2 4 1 -1 ]
  myMUL8 g25 (.A(w15), .B(w17), .Out(w23));   //: @(761, -564) /sz:(170, 138) /sn:0 /p:[ Ti0>0 Ri0>0 Bo0<7 ]
  MYREGISTER18 g29 (.Clk(clk), .in(w18), .out(w22));   //: @(918, -262) /sz:(123, 41) /sn:0 /p:[ Li0>3 Li1>0 Ro0<9 ]
  //: LED g17 (delta) @(1554,417) /sn:0 /w:[ 5 ] /type:3
  //: LED g62 (w22) @(981,-312) /sn:0 /w:[ 7 ] /type:1
  MYREGISTER8 g42 (.in(w20), .Clk(clk), .out(w25));   //: @(173, -371) /sz:(106, 88) /R:3 /sn:0 /p:[ Ti0>0 Ti1>19 Bo0<0 ]
  //: joint g52 (w22) @(1068, -250) /w:[ 1 2 8 -1 ]
  //: joint g63 (w22) @(1068, -291) /w:[ -1 4 6 3 ]
  //: LED g5 (w3) @(568,313) /sn:0 /w:[ 0 ] /type:0
  MYREGISTER18 g14 (.Clk(clk), .in(w12), .out(w16));   //: @(981, 0) /sz:(123, 41) /R:2 /sn:0 /p:[ Ri0>0 Ri1>0 Lo0<0 ]
  //: LED g56 (w16) @(1117,182) /sn:0 /w:[ 5 ] /type:1
  myMUL8 g44 (.A(w25), .B(w25), .Out(w26));   //: @(168, -219) /sz:(170, 138) /sn:0 /p:[ Ti0>5 Ri0>3 Bo0<1 ]
  //: GROUND g47 (w19) @(177,9) /sn:0 /w:[ 0 ]
  MYREGISTER8 g24 (.Clk(clk), .in(c), .out(w17));   //: @(986, -672) /sz:(88, 106) /sn:0 /p:[ Li0>13 Li1>9 Ro0<1 ]
  //: LED g21 (w0) @(989,418) /sn:0 /w:[ 5 ] /type:3
  //: DIP g36 (b) @(254,-724) /sn:0 /w:[ 5 ] /st:3 /dn:1
  MYREGISTER8 g23 (.Clk(clk), .in(a), .out(w15));   //: @(720, -676) /sz:(88, 106) /sn:0 /p:[ Li0>11 Li1>7 Ro0<1 ]
  //: joint g41 (w21) @(714, -343) /w:[ 2 1 4 -1 ]
  //: GROUND g40 (w21) @(664,-320) /sn:0 /w:[ 5 ]
  //: LED g54 (w9) @(1213,397) /sn:0 /w:[ 0 ] /type:0
  //: LED g60 (w23) @(647,-434) /sn:0 /w:[ 9 ] /type:1
  //: LED g70 (c) @(1124,-718) /sn:0 /w:[ 5 ] /type:1
  //: joint g26 (clk) @(667, -586) /w:[ 10 -1 9 12 ]
  MYADDER18 g0 (.A(w8), .B(w16), .Cin(w6), .Cout(w3), .S(w11));   //: @(609, 295) /sz:(164, 142) /sn:0 /p:[ Ti0>5 Ti1>9 Ri0>1 Lo0<1 Bo0<1 ]
  assign w18 = {w23, w21, w21}; //: CONCAT g35  @(793,-353) /sn:0 /w:[ 1 0 0 3 ] /dr:0 /tp:0 /drp:1
  //: joint g45 (w25) @(246, -247) /w:[ 2 1 -1 4 ]
  assign w27 = {w19, w19, w26}; //: CONCAT g46  @(326,-26) /sn:0 /w:[ 1 3 5 0 ] /dr:1 /tp:0 /drp:1
  //: joint g22 (w4) @(1058, 503) /w:[ 2 1 -1 4 ]
  //: LED g66 (b) @(352,-728) /sn:0 /w:[ 3 ] /type:3
  //: joint g12 (w0) @(989, 476) /w:[ 3 4 6 8 ]
  //: joint g18 (delta) @(1554, 475) /w:[ 2 4 1 -1 ]
  //: LED g30 (a) @(768,-735) /sn:0 /w:[ 3 ] /type:3
  //: joint g33 (c) @(962, -682) /w:[ 2 1 -1 8 ]
  MYREGISTER18 g49 (.Clk(clk), .in(w27), .out(w8));   //: @(337, 23) /sz:(41, 123) /R:3 /sn:0 /p:[ Ti0>31 Ti1>0 Bo0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin MYADDER4
module MYADDER4(Cin, A, B, S, Cout);
//: interface  /sz:(145, 40) /bd:[ Ti0>B[3:0](97/145) Ti1>A[3:0](36/145) Ri0>Cin(12/40) Lo0<Cout(12/40) Bo0<S[3:0](71/145) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [3:0] B;    //: /sn:0 {0}(#:32,103)(285,103){1}
//: {2}(286,103)(457,103){3}
//: {4}(458,103)(636,103){5}
//: {6}(637,103)(826,103){7}
//: {8}(827,103)(929,103)(929,95){9}
input [3:0] A;    //: /sn:0 {0}(#:44,57)(241,57){1}
//: {2}(242,57)(411,57){3}
//: {4}(412,57)(590,57){5}
//: {6}(591,57)(773,57){7}
//: {8}(774,57)(932,57){9}
output Cout;    //: /sn:0 {0}(228,208)(162,208)(162,220)(133,220){1}
input Cin;    //: /sn:0 {0}(938,209)(852,209){1}
output [3:0] S;    //: /sn:0 {0}(#:859,332)(951,332)(951,337)(966,337){1}
wire w6;    //: /sn:0 {0}(458,107)(458,138)(466,138)(466,170){1}
wire w7;    //: /sn:0 {0}(320,209)(394,209)(394,208)(399,208){1}
wire w16;    //: /sn:0 {0}(827,107)(827,170){1}
wire w15;    //: /sn:0 {0}(774,61)(774,115)(783,115)(783,170){1}
wire w0;    //: /sn:0 {0}(242,61)(242,115)(251,115)(251,170){1}
wire w3;    //: /sn:0 {0}(807,260)(807,347)(853,347){1}
wire w1;    //: /sn:0 {0}(286,107)(286,115)(295,115)(295,170){1}
wire w8;    //: /sn:0 {0}(624,260)(624,337)(853,337){1}
wire w18;    //: /sn:0 {0}(275,260)(275,317)(853,317){1}
wire w17;    //: /sn:0 {0}(577,208)(569,208){1}
//: {2}(565,208)(527,208)(527,209)(491,209){3}
//: {4}(567,210)(567,217){5}
wire w11;    //: /sn:0 {0}(637,107)(637,115)(644,115)(644,170){1}
wire w10;    //: /sn:0 {0}(591,61)(591,115)(600,115)(600,170){1}
wire w13;    //: /sn:0 {0}(446,260)(446,327)(853,327){1}
wire w5;    //: /sn:0 {0}(412,61)(412,69)(422,69)(422,170){1}
wire w9;    //: /sn:0 {0}(760,208)(725,208)(725,209)(669,209){1}
//: enddecls

  //: IN g4 (Cin) @(940,209) /sn:0 /R:2 /w:[ 0 ]
  assign w0 = A[3]; //: TAP g8 @(242,55) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  FA g3 (.A(w15), .B(w16), .Cin(Cin), .Cout(w9), .S(w3));   //: @(761, 171) /sz:(90, 88) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  assign w11 = B[1]; //: TAP g13 @(637,101) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  FA g2 (.A(w10), .B(w11), .Cin(w9), .Cout(w17), .S(w8));   //: @(578, 171) /sz:(90, 88) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  FA g1 (.A(w5), .B(w6), .Cin(w17), .Cout(w7), .S(w13));   //: @(400, 171) /sz:(90, 88) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>3 Lo0<1 Bo0<0 ]
  assign w6 = B[2]; //: TAP g11 @(458,101) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  assign S = {w18, w13, w8, w3}; //: CONCAT g16  @(858,332) /sn:0 /w:[ 0 1 1 1 1 ] /dr:0 /tp:0 /drp:1
  assign w5 = A[2]; //: TAP g10 @(412,55) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: IN g6 (A) @(42,57) /sn:0 /w:[ 0 ]
  //: IN g7 (B) @(30,103) /sn:0 /w:[ 0 ]
  assign w1 = B[3]; //: TAP g9 @(286,101) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  assign w16 = B[0]; //: TAP g15 @(827,101) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  //: OUT g17 (S) @(963,337) /sn:0 /w:[ 1 ]
  //: OUT g5 (Cout) @(136,220) /sn:0 /R:2 /w:[ 1 ]
  assign w15 = A[0]; //: TAP g14 @(774,55) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  FA g0 (.A(w0), .B(w1), .Cin(w7), .Cout(Cout), .S(w18));   //: @(229, 171) /sz:(90, 88) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<0 ]
  assign w10 = A[1]; //: TAP g12 @(591,55) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  //: joint g18 (w17) @(567, 208) /w:[ 1 -1 2 4 ]

endmodule
//: /netlistEnd

//: /netlistBegin MYADDER2
module MYADDER2(Cout, B, A, S, Cin);
//: interface  /sz:(138, 52) /bd:[ Ti0>B[1:0](90/138) Ti1>A[1:0](33/138) Ri0>Cin(18/52) Lo0<Cout(19/52) Bo0<S[1:0](65/138) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [1:0] B;    //: /sn:0 {0}(#:50,77)(276,77){1}
//: {2}(277,77)(498,77){3}
//: {4}(499,77)(673,77){5}
input [1:0] A;    //: /sn:0 {0}(#:67,46)(235,46){1}
//: {2}(236,46)(447,46){3}
//: {4}(448,46)(650,46){5}
output Cout;    //: /sn:0 {0}(214,205)(153,205)(153,204)(141,204){1}
input Cin;    //: /sn:0 {0}(525,206)(607,206){1}
output [1:0] S;    //: /sn:0 {0}(#:579,303)(609,303)(609,302)(624,302){1}
wire w6;    //: /sn:0 {0}(456,167)(456,58)(448,58)(448,50){1}
wire w4;    //: /sn:0 {0}(480,257)(480,308)(573,308){1}
wire w0;    //: /sn:0 {0}(281,167)(281,89)(277,89)(277,81){1}
wire w3;    //: /sn:0 {0}(306,206)(398,206)(398,205)(433,205){1}
wire w1;    //: /sn:0 {0}(237,167)(237,58)(236,58)(236,50){1}
wire w5;    //: /sn:0 {0}(500,167)(500,89)(499,89)(499,81){1}
wire w9;    //: /sn:0 {0}(261,257)(261,298)(573,298){1}
//: enddecls

  //: OUT g8 (Cout) @(144,204) /sn:0 /R:2 /w:[ 1 ]
  assign w1 = A[1]; //: TAP g4 @(236,44) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  //: IN g3 (B) @(48,77) /sn:0 /w:[ 0 ]
  //: IN g2 (A) @(65,46) /sn:0 /w:[ 0 ]
  FA g1 (.A(w6), .B(w5), .Cin(Cin), .Cout(w3), .S(w4));   //: @(434, 168) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<1 Bo0<0 ]
  //: OUT g11 (S) @(621,302) /sn:0 /w:[ 1 ]
  assign S = {w9, w4}; //: CONCAT g10  @(578,303) /sn:0 /w:[ 0 1 1 ] /dr:0 /tp:0 /drp:1
  assign w6 = A[0]; //: TAP g6 @(448,44) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  //: IN g9 (Cin) @(609,206) /sn:0 /R:2 /w:[ 1 ]
  assign w5 = B[0]; //: TAP g7 @(499,75) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  assign w0 = B[1]; //: TAP g5 @(277,75) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  FA g0 (.A(w1), .B(w0), .Cin(w3), .Cout(Cout), .S(w9));   //: @(215, 168) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<0 Bo0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin latchSR
module latchSR(Y1, R, S, Y);
//: interface  /sz:(101, 105) /bd:[ Li0>S(25/105) Li1>R(80/105) Ri0>Y(81/105) Ro0<Y1(27/105) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input R;    //: /sn:0 {0}(129,308)(266,308)(266,309)(287,309){1}
input S;    //: /sn:0 {0}(146,130)(287,130){1}
output Y1;    //: /sn:0 {0}(521,149)(437,149){1}
//: {2}(433,149)(419,149)(419,148)(406,148){3}
//: {4}(435,151)(435,225)(277,225)(277,268)(287,268){5}
output Y;    //: /sn:0 {0}(536,293)(447,293){1}
//: {2}(445,291)(445,206)(277,206)(277,171)(287,171){3}
//: {4}(443,293)(419,293)(419,286)(406,286){5}
//: enddecls

  //: OUT g4 (Y1) @(518,149) /sn:0 /w:[ 0 ]
  //: IN g3 (R) @(127,308) /sn:0 /w:[ 0 ]
  //: IN g2 (S) @(144,130) /sn:0 /w:[ 0 ]
  myNOR g1 (.in1(Y1), .in2(R), .out(Y));   //: @(288, 239) /sz:(117, 91) /sn:0 /p:[ Li0>5 Li1>1 Ro0<5 ]
  //: joint g6 (Y) @(445, 293) /w:[ 1 2 4 -1 ]
  //: joint g7 (Y1) @(435, 149) /w:[ 1 -1 2 4 ]
  //: OUT g5 (Y) @(533,293) /sn:0 /w:[ 0 ]
  myNOR g0 (.in1(S), .in2(Y), .out(Y1));   //: @(288, 101) /sz:(117, 91) /sn:0 /p:[ Li0>1 Li1>3 Ro0<3 ]

endmodule
//: /netlistEnd

//: /netlistBegin myMUL8
module myMUL8(B, A, Out);
//: interface  /sz:(170, 138) /bd:[ Ti0>A[7:0](78/170) Ri0>B[7:0](69/138) Bo0<Out[15:0](89/170) ] /pd: 0 /pi: 1 /pe: 1 /pp: 1
//: property prot_intf=1
input [7:0] A;    //: {0}(#:-1017,2394)(-976,2394){1}
//: {2}(-975,2394)(-816,2394){3}
//: {4}(-815,2394)(-674,2394){5}
//: {6}(-673,2394)(-539,2394){7}
//: {8}(-538,2394)(-413,2394){9}
//: {10}(-412,2394)(-277,2394){11}
//: {12}(-276,2394)(-143,2394){13}
//: {14}(-142,2394)(-13,2394){15}
//: {16}(-12,2394)(656,2394)(#:656,1997){17}
//: {18}(656,1993)(656,1668){19}
//: {20}(656,1664)(656,1325){21}
//: {22}(656,1321)(656,982){23}
//: {24}(656,978)(656,802)(657,802)(657,627){25}
//: {26}(657,623)(657,463)(664,463)(664,303){27}
//: {28}(666,301)(706,301){29}
//: {30}(662,301)(569,301){31}
//: {32}(568,301)(499,301)(499,300)(432,300){33}
//: {34}(431,300)(371,300)(371,301)(312,301){35}
//: {36}(311,301)(196,301){37}
//: {38}(195,301)(91,301){39}
//: {40}(90,301)(-7,301){41}
//: {42}(-8,301)(-110,301){43}
//: {44}(-111,301)(-212,301){45}
//: {46}(-213,301)(-284,301)(-284,62){47}
//: {48}(-282,60)(-145,60){49}
//: {50}(-144,60)(-40,60){51}
//: {52}(-39,60)(57,60){53}
//: {54}(58,60)(161,60){55}
//: {56}(162,60)(272,60){57}
//: {58}(273,60)(383,60){59}
//: {60}(384,60)(519,60){61}
//: {62}(520,60)(582,60)(582,61)(645,61){63}
//: {64}(646,61)(656,61){65}
//: {66}(-286,60)(#:-330,60){67}
//: {68}(655,625)(479,625){69}
//: {70}(478,625)(350,625){71}
//: {72}(349,625)(240,625){73}
//: {74}(239,625)(134,625){75}
//: {76}(133,625)(30,625){77}
//: {78}(29,625)(-88,625){79}
//: {80}(-89,625)(-207,625){81}
//: {82}(-208,625)(-314,625){83}
//: {84}(-315,625)(-369,625){85}
//: {86}(654,980)(534,980)(534,974)(424,974){87}
//: {88}(423,974)(375,974)(375,980)(336,980){89}
//: {90}(335,980)(228,980){91}
//: {92}(227,980)(119,980){93}
//: {94}(118,980)(-14,980){95}
//: {96}(-15,980)(-143,980){97}
//: {98}(-144,980)(-201,980)(-201,989)(-258,989){99}
//: {100}(-259,989)(-331,989)(-331,980)(-403,980){101}
//: {102}(-404,980)(-482,980){103}
//: {104}(654,1323)(359,1323){105}
//: {106}(358,1323)(230,1323){107}
//: {108}(229,1323)(121,1323){109}
//: {110}(120,1323)(13,1323){111}
//: {112}(12,1323)(-102,1323){113}
//: {114}(-103,1323)(-227,1323){115}
//: {116}(-228,1323)(-343,1323){117}
//: {118}(-344,1323)(-468,1323){119}
//: {120}(-469,1323)(-486,1323){121}
//: {122}(86:654,1666)(343,1666)(343,1668)(254,1668){123}
//: {124}(253,1668)(126,1668){125}
//: {126}(125,1668)(-3,1668){127}
//: {128}(-4,1668)(-128,1668){129}
//: {130}(-129,1668)(-243,1668){131}
//: {132}(-244,1668)(-380,1668){133}
//: {134}(-381,1668)(-513,1668){135}
//: {136}(-514,1668)(-633,1668){137}
//: {138}(-634,1668)(#:-756,1668){139}
//: {140}(654,1995)(103,1995){141}
//: {142}(102,1995)(-29,1995){143}
//: {144}(-30,1995)(-151,1995)(-151,1997)(-161,1997){145}
//: {146}(-162,1997)(-293,1997){147}
//: {148}(-294,1997)(-424,1997){149}
//: {150}(-425,1997)(-541,1997)(-541,1996)(-551,1996){151}
//: {152}(-552,1996)(-689,1996){153}
//: {154}(-690,1996)(-821,1996){155}
//: {156}(-822,1996)(#:-1005,1996){157}
output [15:0] Out;    //: /sn:0 {0}(#:-148,3051)(-148,3095){1}
input [7:0] B;    //: /sn:0 {0}(#:814,50)(814,102){1}
//: {2}(814,103)(814,267){3}
//: {4}(814,268)(814,662){5}
//: {6}(814,663)(814,991){7}
//: {8}(814,992)(814,1352){9}
//: {10}(814,1353)(814,1685){11}
//: {12}(814,1686)(814,2028){13}
//: {14}(814,2029)(814,2433){15}
//: {16}(814,2434)(814,2480){17}
wire w32;    //: /sn:0 {0}(-150,518)(-150,501)(-129,501)(-129,454){1}
wire w270;    //: /sn:0 {0}(-296,2965)(-296,2957)(-1167,2957)(-1167,2653)(-1095,2653){1}
wire w160;    //: /sn:0 {0}(84,2194)(84,2223)(41,2223)(41,2229){1}
wire w96;    //: /sn:0 {0}(569,349)(569,305){1}
wire w73;    //: /sn:0 {0}(-74,932)(-82,932)(-82,933)(-95,933){1}
wire w45;    //: /sn:0 {0}(-99,556)(-100,556)(-100,557)(-125,557){1}
wire w214;    //: /sn:0 {0}(-319,2615)(-319,2587)(-295,2587)(-295,2575){1}
wire w203;    //: /sn:0 {0}(-821,2089)(-821,2000){1}
wire w166;    //: /sn:0 {0}(-446,1576)(-473,1576){1}
wire w134;    //: /sn:0 {0}(-344,1378)(-344,1335)(-343,1335)(-343,1327){1}
wire w122;    //: /sn:0 {0}(-122,1222)(-143,1222)(-143,1223)(-158,1223){1}
wire w220;    //: /sn:0 {0}(-537,2470)(-537,2406)(-538,2406)(-538,2398){1}
wire w141;    //: /sn:0 {0}(154,1580)(139,1580)(139,1579)(128,1579){1}
wire w14;    //: /sn:0 {0}(143,232)(143,301)(126,301)(126,504)(144,504)(144,517){1}
wire w218;    //: /sn:0 {0}(-363,2615)(-363,2485)(-359,2485)(-359,2327){1}
wire w56;    //: /sn:0 {0}(-7,894)(-7,852)(12,852)(12,827){1}
wire w16;    //: /sn:0 {0}(429,517)(429,500)(414,500)(414,454){1}
wire w179;    //: /sn:0 {0}(-98,1898)(-121,1898)(-121,1897)(-136,1897){1}
wire w81;    //: /sn:0 {0}(-270,1025)(-270,1014)(-258,1014)(-258,993){1}
wire w89;    //: /sn:0 {0}(-351,1184)(-351,1000)(-382,1000)(-382,984){1}
wire w4;    //: /sn:0 {0}(-352,722)(-352,663)(-218,663){1}
//: {2}(-214,663)(-116,663){3}
//: {4}(-112,663)(-9,663){5}
//: {6}(-5,663)(95,663){7}
//: {8}(99,663)(202,663){9}
//: {10}(206,663)(311,663){11}
//: {12}(315,663)(439,663){13}
//: {14}(443,663)(809,663){15}
//: {16}(441,665)(441,691)(441,691)(441,722){17}
//: {18}(313,665)(313,692)(313,692)(313,722){19}
//: {20}(204,665)(204,722){21}
//: {22}(97,665)(97,692)(97,692)(97,722){23}
//: {24}(-7,665)(-7,693)(-7,693)(-7,722){25}
//: {26}(-114,665)(-114,694)(-126,694)(-126,722){27}
//: {28}(-216,665)(-216,690)(-245,690)(-245,717){29}
wire w19;    //: /sn:0 {0}(366,232)(366,482)(385,482)(385,517){1}
wire w266;    //: /sn:0 {0}(-276,2965)(-276,2949)(-906,2949)(-906,2705){1}
wire w250;    //: /sn:0 {0}(-560,2654)(-532,2654)(-532,2653)(-514,2653){1}
wire w195;    //: /sn:0 {0}(-511,2237)(-511,1994)(-435,1994)(-435,1944){1}
wire w38;    //: /sn:0 {0}(354,933)(365,933)(365,918)(424,918){1}
wire w182;    //: /sn:0 {0}(-205,2238)(-205,2209)(-180,2209)(-180,2194){1}
wire w180;    //: /sn:0 {0}(-119,2237)(-119,2000)(-51,2000)(-51,1950){1}
wire w152;    //: /sn:0 {0}(-75,1860)(-75,1643)(-34,1643)(-34,1628){1}
wire w183;    //: /sn:0 {0}(12,2271)(-44,2271)(-44,2276)(-50,2276){1}
wire w181;    //: /sn:0 {0}(-228,1896)(-247,1896){1}
wire w194;    //: /sn:0 {0}(-482,1892)(-512,1892)(-512,1896)(-516,1896){1}
wire w3;    //: /sn:0 {0}(647,127)(647,96)(646,96)(646,65){1}
wire w151;    //: /sn:0 {0}(-81,1576)(-94,1576)(-94,1577)(-109,1577){1}
wire w0;    //: /sn:0 {0}(460,827)(460,842)(453,842)(453,876){1}
wire w128;    //: /sn:0 {0}(-178,1538)(-178,1289)(-203,1289)(-203,1274){1}
wire w127;    //: /sn:0 {0}(-250,1222)(-267,1222)(-267,1223)(-282,1223){1}
wire w240;    //: /sn:0 {0}(-252,2653)(-270,2653)(-270,2654)(-294,2654){1}
wire w233;    //: /sn:0 {0}(-767,2615)(-767,2341)(-760,2341)(-760,2326){1}
wire w120;    //: /sn:0 {0}(-35,2965)(-35,2937)(310,2937)(310,1641)(328,1641)(328,1626){1}
wire w133;    //: /sn:0 {0}(-306,1539)(-306,1289)(-327,1289)(-327,1274){1}
wire w168;    //: /sn:0 {0}(-541,1857)(-541,1832)(-530,1832)(-530,1823){1}
wire w171;    //: /sn:0 {0}(-565,1575)(-716,1575)(-716,1856){1}
wire w111;    //: /sn:0 {0}(122,1373)(122,1335)(121,1335)(121,1327){1}
wire w104;    //: /sn:0 {0}(339,1477)(339,1487)(302,1487)(302,1538){1}
wire w204;    //: /sn:0 {0}(-739,1894)(-939,1894)(-939,2236){1}
wire w75;    //: /sn:0 {0}(-55,1184)(-55,1144)(-32,1144)(-32,1130){1}
wire w237;    //: /sn:0 {0}(-962,2274)(-1072,2274)(-1072,2615){1}
wire w209;    //: /sn:0 {0}(-185,2615)(-185,2587)(-161,2587)(-161,2575){1}
wire w119;    //: /sn:0 {0}(-14,1538)(-14,1494)(-4,1494)(-4,1479){1}
wire w67;    //: /sn:0 {0}(59,127)(59,105)(59,105)(59,68)(58,68)(58,64){1}
wire w54;    //: /sn:0 {0}(-406,894)(-406,546)(-355,546){1}
wire w215;    //: /sn:0 {0}(-412,2470)(-412,2398){1}
wire w176;    //: /sn:0 {0}(-75,2237)(-75,2209)(-48,2209)(-48,2194){1}
wire w90;    //: /sn:0 {0}(-428,1184)(-428,1148)(-410,1148)(-410,1130){1}
wire w156;    //: /sn:0 {0}(-201,1576)(-222,1576)(-222,1578)(-237,1578){1}
wire w167;    //: /sn:0 {0}(-459,1854)(-459,1640)(-399,1640)(-399,1628){1}
wire w41;    //: /sn:0 {0}(-212,349)(-212,305){1}
wire w36;    //: /sn:0 {0}(415,1130)(415,1147)(397,1147)(397,1178){1}
wire w174;    //: /sn:0 {0}(33,1901)(9,1901)(9,1899)(-6,1899){1}
wire w124;    //: /sn:0 {0}(-134,1538)(-134,1496)(-121,1496)(-121,1481){1}
wire w23;    //: /sn:0 {0}(-163,232)(-163,484)(-194,484)(-194,518){1}
wire w20;    //: /sn:0 {0}(-76,518)(-76,486)(-57,486)(-57,232){1}
wire w225;    //: /sn:0 {0}(-671,2470)(-671,2406)(-673,2406)(-673,2398){1}
wire w108;    //: /sn:0 {0}(363,1538)(363,1319)(292,1319)(292,1274){1}
wire w82;    //: /sn:0 {0}(273,127)(273,106)(273,106)(273,64){1}
wire w223;    //: /sn:0 {0}(-491,2615)(-491,2485)(-487,2485)(-487,2327){1}
wire w126;    //: /sn:0 {0}(235,1835)(235,1854)(224,1854)(224,1840)(191,1840)(191,1864){1}
wire w158;    //: /sn:0 {0}(-272,1857)(-272,1838)(-262,1838)(-262,1823){1}
wire w74;    //: /sn:0 {0}(34,1184)(34,997)(-27,997)(-27,984){1}
wire w125;    //: /sn:0 {0}(-227,1184)(-227,999)(-264,999)(-264,984){1}
wire w91;    //: /sn:0 {0}(242,722)(242,637)(240,637)(240,629){1}
wire w35;    //: /sn:0 {0}(121,555)(112,555)(112,556)(110,556){1}
wire w8;    //: /sn:0 {0}(-231,454)(-231,464)(-265,464)(-265,504){1}
wire w103;    //: /sn:0 {0}(-25,2965)(-25,2941)(423,2941)(423,1266){1}
wire w192;    //: /sn:0 {0}(-31,2575)(-31,2585)(-87,2585)(-87,2605){1}
wire w163;    //: /sn:0 {0}(-415,1854)(-415,1835)(-399,1835)(-399,1823){1}
wire w101;    //: /sn:0 {0}(358,1372)(358,1342)(359,1342)(359,1327){1}
wire w238;    //: /sn:0 {0}(-915,2326)(-915,2605)(-930,2605)(-930,2615){1}
wire w71;    //: /sn:0 {0}(-13,1025)(-13,992)(-14,992)(-14,984){1}
wire w144;    //: /sn:0 {0}(-859,2089)(-859,2029)(-730,2029){1}
//: {2}(-726,2029)(-712,2029)(-712,2029)(-591,2029){3}
//: {4}(-587,2029)(-464,2029){5}
//: {6}(-460,2029)(-332,2029){7}
//: {8}(-328,2029)(-201,2029){9}
//: {10}(-197,2029)(-69,2029){11}
//: {12}(-65,2029)(63,2029){13}
//: {14}(67,2029)(809,2029){15}
//: {16}(65,2031)(65,2089){17}
//: {18}(-67,2031)(-67,2089){19}
//: {20}(-199,2031)(-199,2089){21}
//: {22}(-330,2031)(-330,2060)(-329,2060)(-329,2089){23}
//: {24}(-462,2031)(-462,2089){25}
//: {26}(-589,2031)(-589,2089){27}
//: {28}(-728,2031)(-728,2089){29}
wire w22;    //: /sn:0 {0}(-5,2965)(-5,2952)(546,2952)(546,600){1}
wire w265;    //: /sn:0 {0}(-953,2653)(-975,2653)(-975,2654)(-1003,2654){1}
wire w17;    //: /sn:0 {0}(40,232)(40,313)(41,313)(41,517){1}
wire w117;    //: /sn:0 {0}(11,1222)(-6,1222)(-6,1223)(-30,1223){1}
wire w53;    //: /sn:0 {0}(309,984)(309,994)(458,994)(458,1178){1}
wire w172;    //: /sn:0 {0}(-585,1857)(-585,1636)(-518,1636)(-518,1627){1}
wire w255;    //: /sn:0 {0}(-652,2653)(-686,2653)(-686,2654)(-698,2654){1}
wire w228;    //: /sn:0 {0}(-629,2615)(-629,2485)(-625,2485)(-625,2326){1}
wire w12;    //: /sn:0 {0}(91,305)(91,313)(92,313)(92,349){1}
wire w44;    //: /sn:0 {0}(312,1184)(312,1142)(317,1142)(317,1130){1}
wire w2;    //: /sn:0 {0}(628,232)(628,2958)(5,2958)(5,2965){1}
wire w113;    //: /sn:0 {0}(186,1274)(186,1313)(161,1313)(161,1532)(177,1532)(177,1542){1}
wire [7:0] w226;    //: /sn:0 {0}(-143,3045)(-143,2986)(#:-30,2986)(#:-30,2971){1}
wire w115;    //: /sn:0 {0}(246,1581)(270,1581)(270,1580)(273,1580){1}
wire w77;    //: /sn:0 {0}(162,127)(162,106)(162,106)(162,64){1}
wire w83;    //: /sn:0 {0}(-337,933)(-327,933)(-327,932)(-311,932){1}
wire w200;    //: /sn:0 {0}(-649,2236)(-649,1997)(-561,1997)(-561,1947){1}
wire w78;    //: /sn:0 {0}(-187,932)(-211,932)(-211,933)(-219,933){1}
wire w224;    //: /sn:0 {0}(-585,2615)(-585,2590)(-556,2590)(-556,2575){1}
wire w10;    //: /sn:0 {0}(550,454)(550,467)(520,467)(520,512){1}
wire w27;    //: /sn:0 {0}(362,555)(350,555)(350,556)(332,556){1}
wire w190;    //: /sn:0 {0}(-383,2237)(-383,1997)(-292,1997)(-292,1947){1}
wire w246;    //: /sn:0 {0}(-236,2965)(-236,2908)(-339,2908)(-339,2705){1}
wire w138;    //: /sn:0 {0}(-448,1274)(-448,1311)(-423,1311)(-423,1538){1}
wire w86;    //: /sn:0 {0}(-391,1025)(-391,992)(-403,992)(-403,984){1}
wire w188;    //: /sn:0 {0}(-424,2089)(-424,2001){1}
wire w95;    //: /sn:0 {0}(479,629)(479,722){1}
wire w52;    //: /sn:0 {0}(119,1025)(119,984){1}
wire w80;    //: /sn:0 {0}(-183,1184)(-183,1144)(-162,1144)(-162,1130){1}
wire w29;    //: /sn:0 {0}(385,127)(385,106)(385,106)(385,68)(384,68)(384,64){1}
wire w187;    //: /sn:0 {0}(-55,2965)(-55,2926)(67,2926)(67,2317){1}
wire w178;    //: /sn:0 {0}(-161,2089)(-161,2001){1}
wire w155;    //: /sn:0 {0}(-45,2965)(-45,2932)(217,2932)(217,1952){1}
wire w142;    //: /sn:0 {0}(201,1632)(201,1639)(252,1639)(252,1864){1}
wire w147;    //: /sn:0 {0}(56,1863)(56,1645)(83,1645)(83,1630){1}
wire w42;    //: /sn:0 {0}(-15,2965)(-15,2945)(479,2945)(479,964){1}
wire w50;    //: /sn:0 {0}(-217,556)(-287,556)(-287,521)(-276,521)(-276,491)(-311,491)(-311,479)(-326,479)(-326,504){1}
wire w6;    //: /sn:0 {0}(519,127)(519,68)(520,68)(520,64){1}
wire w93;    //: /sn:0 {0}(350,629)(350,637)(351,637)(351,722){1}
wire w7;    //: /sn:0 {0}(-250,349)(-250,268)(-150,268){1}
//: {2}(-146,268)(-47,268){3}
//: {4}(-43,268)(52,268){5}
//: {6}(56,268)(156,268){7}
//: {8}(160,268)(272,268){9}
//: {10}(276,268)(393,268){11}
//: {12}(397,268)(529,268){13}
//: {14}(533,268)(809,268){15}
//: {16}(531,270)(531,311)(531,311)(531,349){17}
//: {18}(395,270)(395,310)(395,310)(395,349){19}
//: {20}(274,270)(274,310)(274,310)(274,349){21}
//: {22}(158,270)(158,310)(158,310)(158,349){23}
//: {24}(54,270)(54,309)(54,309)(54,349){25}
//: {26}(-45,270)(-45,309)(-45,309)(-45,349){27}
//: {28}(-148,270)(-148,308)(-148,308)(-148,349){29}
wire w60;    //: /sn:0 {0}(262,932)(244,932){1}
wire w99;    //: /sn:0 {0}(336,1025)(336,984){1}
wire w61;    //: /sn:0 {0}(152,931)(141,931)(141,933)(123,933){1}
wire w46;    //: /sn:0 {0}(-52,608)(-52,766)(-51,766)(-51,894){1}
wire w175;    //: /sn:0 {0}(80,1953)(80,2040)(147,2040)(147,2218)(102,2218)(102,2229){1}
wire w112;    //: /sn:0 {0}(139,1222)(124,1222)(124,1223)(103,1223){1}
wire w135;    //: /sn:0 {0}(-363,1483)(-363,1523)(-379,1523)(-379,1538){1}
wire w153;    //: /sn:0 {0}(-161,1858)(-161,1833)(-146,1833)(-146,1823){1}
wire w216;    //: /sn:0 {0}(-160,2654)(-140,2654)(-140,2647)(-116,2647){1}
wire w15;    //: /sn:0 {0}(-88,629)(-88,722){1}
wire w207;    //: /sn:0 {0}(-142,2275)(-165,2275)(-165,2277)(-180,2277){1}
wire w213;    //: /sn:0 {0}(-229,2615)(-229,2485)(-225,2485)(-225,2328){1}
wire w239;    //: /sn:0 {0}(-1028,2615)(-1028,2591)(-993,2591)(-993,2575){1}
wire w106;    //: /sn:0 {0}(232,1373)(232,1335)(230,1335)(230,1327){1}
wire w51;    //: /sn:0 {0}(-170,608)(-170,913)(-179,913)(-179,884)(-164,884)(-164,894){1}
wire w69;    //: /sn:0 {0}(162,1184)(162,995)(78,995)(78,984){1}
wire w129;    //: /sn:0 {0}(-226,1379)(-226,1335)(-227,1335)(-227,1327){1}
wire w109;    //: /sn:0 {0}(213,1478)(213,1527)(221,1527)(221,1542){1}
wire w229;    //: /sn:0 {0}(-723,2615)(-723,2590)(-690,2590)(-690,2575){1}
wire w114;    //: /sn:0 {0}(103,1540)(103,1478){1}
wire w97;    //: /sn:0 {0}(135,722)(135,637)(134,637)(134,629){1}
wire w271;    //: /sn:0 {0}(-286,2965)(-286,2954)(-1048,2954)(-1048,2705){1}
wire w177;    //: /sn:0 {0}(-1012,2470)(-1012,2434)(-855,2434){1}
//: {2}(-851,2434)(-711,2434){3}
//: {4}(-707,2434)(-577,2434){5}
//: {6}(-573,2434)(-452,2434){7}
//: {8}(-448,2434)(-316,2434){9}
//: {10}(-312,2434)(-182,2434){11}
//: {12}(-178,2434)(-52,2434){13}
//: {14}(-48,2434)(809,2434){15}
//: {16}(-50,2436)(-50,2470){17}
//: {18}(-180,2436)(-180,2470){19}
//: {20}(-314,2436)(-314,2470){21}
//: {22}(-450,2436)(-450,2470){23}
//: {24}(-575,2436)(-575,2470){25}
//: {26}(-709,2436)(-709,2470){27}
//: {28}(-853,2436)(-853,2470){29}
wire w66;    //: /sn:0 {0}(65,607)(65,884)(54,884)(54,894){1}
wire w37;    //: /sn:0 {0}(409,607)(409,852)(514,852)(514,876){1}
wire w261;    //: /sn:0 {0}(-743,2705)(-743,2937)(-266,2937)(-266,2965){1}
wire w64;    //: /sn:0 {0}(98,894)(98,838)(116,838)(116,827){1}
wire w245;    //: /sn:0 {0}(-386,2653)(-406,2653)(-406,2654)(-422,2654){1}
wire w234;    //: /sn:0 {0}(-886,2615)(-886,2590)(-834,2590)(-834,2575){1}
wire w34;    //: /sn:0 {0}(285,894)(285,750)(287,750)(287,607){1}
wire w63;    //: /sn:0 {0}(268,1184)(268,984)(199,984)(199,983){1}
wire w159;    //: /sn:0 {0}(-380,1718)(-380,1672){1}
wire w102;    //: /sn:0 {0}(368,1220)(350,1220)(350,1223)(337,1223){1}
wire w43;    //: /sn:0 {0}(329,894)(329,873)(332,873)(332,827){1}
wire w87;    //: /sn:0 {0}(228,984)(228,1025){1}
wire w157;    //: /sn:0 {0}(-205,1858)(-205,1643)(-154,1643)(-154,1628){1}
wire w21;    //: /sn:0 {0}(-144,127)(-144,108)(-144,108)(-144,64){1}
wire w76;    //: /sn:0 {0}(-143,1025)(-143,984){1}
wire w199;    //: /sn:0 {0}(-608,1895)(-647,1895){1}
wire w170;    //: /sn:0 {0}(-29,2089)(-29,1999){1}
wire w58;    //: /sn:0 {0}(175,893)(175,628)(168,628)(168,607){1}
wire w230;    //: /sn:0 {0}(-815,2470)(-815,2398){1}
wire w31;    //: /sn:0 {0}(-429,1025)(-429,992)(-310,992){1}
//: {2}(-306,992)(-183,992){3}
//: {4}(-179,992)(-53,992){5}
//: {6}(-49,992)(79,992){7}
//: {8}(83,992)(188,992){9}
//: {10}(192,992)(296,992){11}
//: {12}(300,992)(393,992){13}
//: {14}(397,992)(809,992){15}
//: {16}(395,994)(395,1009)(396,1009)(396,1025){17}
//: {18}(298,994)(298,1025){19}
//: {20}(190,994)(190,1025){21}
//: {22}(81,994)(81,1025){23}
//: {24}(-51,994)(-51,1025){25}
//: {26}(-181,994)(-181,1025){27}
//: {28}(-308,994)(-308,1025){29}
wire w100;    //: /sn:0 {0}(434,1025)(434,986)(424,986)(424,978){1}
wire w28;    //: /sn:0 {0}(73,454)(73,501)(85,501)(85,517){1}
wire w130;    //: /sn:0 {0}(-262,1539)(-262,1499)(-245,1499)(-245,1484){1}
wire w169;    //: /sn:0 {0}(-633,1718)(-633,1699)(-633,1699)(-633,1672){1}
wire w24;    //: /sn:0 {0}(293,454)(293,485)(307,485)(307,517){1}
wire w251;    //: /sn:0 {0}(-246,2965)(-246,2918)(-467,2918)(-467,2705){1}
wire w132;    //: /sn:0 {0}(-374,1222)(-394,1222)(-394,1223)(-403,1223){1}
wire w184;    //: /sn:0 {0}(-291,2089)(-291,2044)(-293,2044)(-293,2001){1}
wire w260;    //: /sn:0 {0}(-790,2653)(-845,2653)(-845,2654)(-861,2654){1}
wire w256;    //: /sn:0 {0}(-256,2965)(-256,2927)(-605,2927)(-605,2705){1}
wire w1;    //: /sn:0 {0}(809,103)(611,103){1}
//: {2}(607,103)(483,103){3}
//: {4}(479,103)(349,103){5}
//: {6}(345,103)(237,103){7}
//: {8}(233,103)(126,103){9}
//: {10}(122,103)(23,103){11}
//: {12}(19,103)(-74,103){13}
//: {14}(-78,103)(-182,103)(-182,127){15}
//: {16}(-76,105)(-76,115)(-76,115)(-76,127){17}
//: {18}(21,105)(21,115)(21,115)(21,127){19}
//: {20}(124,105)(124,115)(124,115)(124,127){21}
//: {22}(235,105)(235,115)(235,115)(235,127){23}
//: {24}(347,105)(347,115)(347,115)(347,127){25}
//: {26}(481,105)(481,127){27}
//: {28}(609,105)(609,115)(609,115)(609,127){29}
wire w161;    //: /sn:0 {0}(-329,1577)(-354,1577){1}
wire w235;    //: /sn:0 {0}(-974,2470)(-974,2406)(-975,2406)(-975,2398){1}
wire w140;    //: /sn:0 {0}(-488,1482)(-488,1522)(-498,1522)(-498,1537){1}
wire w196;    //: /sn:0 {0}(-605,2236)(-605,2209)(-570,2209)(-570,2194){1}
wire w221;    //: /sn:0 {0}(-65,2965)(-65,2940)(-61,2940)(-61,2693){1}
wire w241;    //: /sn:0 {0}(-226,2965)(-226,2869)(-205,2869)(-205,2705){1}
wire w25;    //: /sn:0 {0}(-314,629)(-314,722){1}
wire [7:0] w253;    //: /sn:0 {0}(-153,3045)(-153,2986)(#:-261,2986)(#:-261,2971){1}
wire w154;    //: /sn:0 {0}(-243,1718)(-243,1672){1}
wire w205;    //: /sn:0 {0}(-784,2236)(-784,1996)(-692,1996)(-692,1946){1}
wire w65;    //: /sn:0 {0}(-362,894)(-362,841)(-333,841)(-333,827){1}
wire w210;    //: /sn:0 {0}(-276,2470)(-276,2398){1}
wire w98;    //: /sn:0 {0}(-507,1377)(-507,1353)(-384,1353){1}
//: {2}(-380,1353)(-266,1353){3}
//: {4}(-262,1353)(-142,1353){5}
//: {6}(-138,1353)(-25,1353){7}
//: {8}(-21,1353)(82,1353){9}
//: {10}(86,1353)(192,1353){11}
//: {12}(196,1353)(317,1353){13}
//: {14}(321,1353)(809,1353){15}
//: {16}(319,1355)(319,1363)(320,1363)(320,1372){17}
//: {18}(194,1355)(194,1373){19}
//: {20}(84,1355)(84,1373){21}
//: {22}(-23,1355)(-23,1374){23}
//: {24}(-140,1355)(-140,1376){25}
//: {26}(-264,1355)(-264,1379){27}
//: {28}(-382,1355)(-382,1378){29}
wire w116;    //: /sn:0 {0}(15,1374)(15,1335)(13,1335)(13,1327){1}
wire w227;    //: /sn:0 {0}(-672,2274)(-707,2274)(-707,2275)(-715,2275){1}
wire w121;    //: /sn:0 {0}(-102,1376)(-102,1327){1}
wire w92;    //: /sn:0 {0}(312,349)(312,305){1}
wire w40;    //: /sn:0 {0}(18,555)(14,555)(14,557)(-7,557){1}
wire w118;    //: /sn:0 {0}(58,1274)(58,1530)(59,1530)(59,1540){1}
wire w18;    //: /sn:0 {0}(-207,629)(-207,717){1}
wire w212;    //: /sn:0 {0}(-272,2276)(-314,2276){1}
wire w162;    //: /sn:0 {0}(-316,1857)(-316,1644)(-282,1644)(-282,1629){1}
wire w30;    //: /sn:0 {0}(-32,518)(-32,502)(-26,502)(-26,454){1}
wire w217;    //: /sn:0 {0}(-406,2275)(-432,2275)(-432,2276)(-442,2276){1}
wire w164;    //: /sn:0 {0}(-511,1718)(-511,1680)(-513,1680)(-513,1672){1}
wire w68;    //: /sn:0 {0}(31,932)(28,932)(28,933)(18,933){1}
wire w146;    //: /sn:0 {0}(36,1578)(24,1578)(24,1577)(11,1577){1}
wire w149;    //: /sn:0 {0}(125,1902)(154,1902)(154,1906)(162,1906){1}
wire w222;    //: /sn:0 {0}(-534,2275)(-580,2275){1}
wire w198;    //: /sn:0 {0}(-690,2089)(-690,2044)(-689,2044)(-689,2000){1}
wire w165;    //: /sn:0 {0}(-12,2470)(-12,2398){1}
wire w123;    //: /sn:0 {0}(-58,1538)(-58,1289)(-75,1289)(-75,1274){1}
wire w59;    //: /sn:0 {0}(-120,894)(-120,836)(-107,836)(-107,827){1}
wire w62;    //: /sn:0 {0}(-244,894)(-244,830)(-226,830)(-226,822){1}
wire w85;    //: /sn:0 {0}(-307,1184)(-307,1146)(-289,1146)(-289,1130){1}
wire w185;    //: /sn:0 {0}(-249,2238)(-249,1998)(-181,1998)(-181,1948){1}
wire w136;    //: /sn:0 {0}(-671,1718)(-671,1686)(-551,1686){1}
//: {2}(-547,1686)(-420,1686){3}
//: {4}(-416,1686)(-283,1686){5}
//: {6}(-279,1686)(-171,1686){7}
//: {8}(-167,1686)(-43,1686){9}
//: {10}(-39,1686)(86,1686){11}
//: {12}(90,1686)(213,1686){13}
//: {14}(217,1686)(809,1686){15}
//: {16}(215,1688)(215,1700)(216,1700)(216,1730){17}
//: {18}(88,1688)(88,1694)(88,1694)(88,1718){19}
//: {20}(-41,1688)(-41,1704)(-41,1704)(-41,1718){21}
//: {22}(-169,1688)(-169,1698)(-165,1698)(-165,1718){23}
//: {24}(-281,1688)(-281,1718){25}
//: {26}(-418,1688)(-418,1718){27}
//: {28}(-549,1688)(-549,1718){29}
wire w173;    //: /sn:0 {0}(-652,1823)(-652,1841)(-672,1841)(-672,1856){1}
wire w57;    //: /sn:0 {0}(223,827)(223,849)(219,849)(219,893){1}
wire w49;    //: /sn:0 {0}(209,1130)(209,1169)(206,1169)(206,1184){1}
wire w139;    //: /sn:0 {0}(-469,1377)(-469,1335)(-468,1335)(-468,1327){1}
wire w197;    //: /sn:0 {0}(-142,2470)(-142,2398){1}
wire w11;    //: /sn:0 {0}(263,517)(263,506)(234,506)(234,305)(254,305)(254,232){1}
wire w137;    //: /sn:0 {0}(-495,1222)(-542,1222)(-542,1537){1}
wire w148;    //: /sn:0 {0}(-31,1860)(-31,1838)(-22,1838)(-22,1823){1}
wire w105;    //: /sn:0 {0}(254,1730)(254,1672){1}
wire w150;    //: /sn:0 {0}(-127,1718)(-127,1679)(-128,1679)(-128,1672){1}
wire w70;    //: /sn:0 {0}(78,1184)(78,1143)(100,1143)(100,1130){1}
wire w110;    //: /sn:0 {0}(-3,1672)(-3,1718){1}
wire w189;    //: /sn:0 {0}(-339,1895)(-375,1895)(-375,1893)(-390,1893){1}
wire w193;    //: /sn:0 {0}(-551,2089)(-551,2000){1}
wire w186;    //: /sn:0 {0}(-339,2237)(-339,2210)(-310,2210)(-310,2194){1}
wire w206;    //: /sn:0 {0}(-895,2236)(-895,2202)(-840,2202)(-840,2194){1}
wire w72;    //: /sn:0 {0}(30,629)(30,637)(31,637)(31,722){1}
wire w94;    //: /sn:0 {0}(433,349)(433,324)(432,324)(432,304){1}
wire w13;    //: /sn:0 {0}(500,232)(500,482)(581,482)(581,512){1}
wire w88;    //: /sn:0 {0}(-429,932)(-472,932)(-472,1184){1}
wire w33;    //: /sn:0 {0}(213,556)(229,556)(229,555)(240,555){1}
wire w191;    //: /sn:0 {0}(-467,2237)(-467,2209)(-443,2209)(-443,2194){1}
wire w5;    //: /sn:0 {0}(454,556)(474,556)(474,554)(491,554){1}
wire w48;    //: /sn:0 {0}(-7,305)(-7,349){1}
wire w208;    //: /sn:0 {0}(-95,2327)(-95,2465)(-19,2465)(-19,2592)(-26,2592)(-26,2605){1}
wire w143;    //: /sn:0 {0}(100,1863)(100,1838)(107,1838)(107,1823){1}
wire w107;    //: /sn:0 {0}(245,1222)(241,1222)(241,1223)(231,1223){1}
wire w131;    //: /sn:0 {0}(126,1718)(126,1672){1}
wire w47;    //: /sn:0 {0}(-38,127)(-38,107)(-38,107)(-38,68)(-39,68)(-39,64){1}
wire w219;    //: /sn:0 {0}(-447,2615)(-447,2589)(-431,2589)(-431,2575){1}
wire w9;    //: /sn:0 {0}(196,305)(196,349){1}
wire w79;    //: /sn:0 {0}(-99,1184)(-99,993)(-140,993)(-140,984){1}
wire w145;    //: /sn:0 {0}(103,2089)(103,1999){1}
wire w55;    //: /sn:0 {0}(-288,894)(-288,716)(-300,716)(-300,592){1}
wire w39;    //: /sn:0 {0}(-110,305)(-110,349){1}
wire w201;    //: /sn:0 {0}(-740,2236)(-740,2209)(-709,2209)(-709,2194){1}
wire w232;    //: /sn:0 {0}(-807,2274)(-855,2274)(-855,2275)(-870,2275){1}
wire w26;    //: /sn:0 {0}(188,517)(188,499)(177,499)(177,454){1}
//: enddecls

  myAND2 g165 (.B(w136), .A(w159), .Out(w163));   //: @(-437, 1719) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>27 Ti1>0 Bo0<1 ]
  myAND2 g8 (.B(w1), .A(w67), .Out(w17));   //: @(2, 128) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>19 Ti1>0 Bo0<0 ]
  assign w134 = A[6]; //: TAP g140 @(-343,1321) /sn:0 /R:1 /w:[ 1 118 117 ] /ss:1
  FA g55 (.A(w20), .B(w30), .Cin(w40), .Cout(w45), .S(w46));   //: @(-98, 519) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g37 (w7) @(54, 268) /w:[ 6 -1 5 24 ]
  assign w67 = A[5]; //: TAP g13 @(58,58) /sn:0 /R:1 /w:[ 1 53 54 ] /ss:1
  assign w129 = A[5]; //: TAP g139 @(-227,1321) /sn:0 /R:1 /w:[ 1 116 115 ] /ss:1
  assign w99 = A[1]; //: TAP g111 @(336,978) /sn:0 /R:1 /w:[ 1 90 89 ] /ss:1
  FA g218 (.A(w185), .B(w182), .Cin(w207), .Cout(w212), .S(w213));   //: @(-271, 2239) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  //: joint g176 (w136) @(-549, 1686) /w:[ 2 -1 1 28 ]
  //: IN g1 (B) @(814,48) /sn:0 /R:3 /w:[ 0 ]
  assign w21 = A[7]; //: TAP g11 @(-144,58) /sn:0 /R:1 /w:[ 1 49 50 ] /ss:1
  myAND2 g130 (.A(w121), .B(w98), .Out(w124));   //: @(-159, 1377) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>0 Ti1>25 Bo0<1 ]
  MyHA g50 (.B(w10), .A(w13), .cout(w5), .S(w22));   //: @(492, 513) /sz:(107, 86) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<1 ]
  assign w197 = A[1]; //: TAP g254 @(-142,2392) /sn:0 /R:1 /w:[ 1 13 14 ] /ss:1
  FA g223 (.A(w204), .B(w206), .Cin(w232), .Cout(w237), .S(w238));   //: @(-961, 2237) /sz:(90, 88) /sn:0 /p:[ Ti0>1 Ti1>0 Ri0>1 Lo0<0 Bo0<0 ]
  assign w145 = A[0]; //: TAP g197 @(103,1993) /sn:0 /R:1 /w:[ 1 142 141 ] /ss:1
  myAND2 g132 (.A(w134), .B(w98), .Out(w135));   //: @(-401, 1379) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>0 Ti1>29 Bo0<0 ]
  assign w52 = A[3]; //: TAP g113 @(119,978) /sn:0 /R:1 /w:[ 1 94 93 ] /ss:1
  //: joint g19 (w1) @(609, 103) /w:[ 1 -1 2 28 ]
  MyHA g150 (.B(w104), .A(w108), .cout(w115), .S(w120));   //: @(274, 1539) /sz:(107, 86) /sn:0 /p:[ Ti0>1 Ti1>0 Lo0<1 Bo0<1 ]
  //: joint g146 (w98) @(-23, 1353) /w:[ 8 -1 7 22 ]
  assign w76 = A[5]; //: TAP g115 @(-143,978) /sn:0 /R:1 /w:[ 1 98 97 ] /ss:1
  //: joint g38 (w7) @(-45, 268) /w:[ 4 -1 3 26 ]
  //: joint g75 (A) @(664, 301) /w:[ 28 -1 30 27 ]
  myAND2 g227 (.B(w177), .A(w210), .Out(w214));   //: @(-333, 2471) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>21 Ti1>0 Bo0<1 ]
  assign w136 = B[5]; //: TAP g169 @(812,1686) /sn:0 /R:2 /w:[ 15 12 11 ] /ss:0
  myAND2 g160 (.B(w136), .A(w105), .Out(w126));   //: @(197, 1731) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>17 Ti1>0 Bo0<0 ]
  assign w106 = A[1]; //: TAP g135 @(230,1321) /sn:0 /R:1 /w:[ 1 108 107 ] /ss:1
  myAND2 g31 (.B(w7), .A(w39), .Out(w32));   //: @(-167, 350) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>29 Ti1>1 Bo0<1 ]
  //: joint g20 (w1) @(481, 103) /w:[ 3 -1 4 26 ]
  myAND2 g230 (.B(w177), .A(w225), .Out(w229));   //: @(-728, 2471) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>27 Ti1>0 Bo0<1 ]
  FA g124 (.A(w89), .B(w85), .Cin(w127), .Cout(w132), .S(w133));   //: @(-373, 1185) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  //: joint g68 (w4) @(313, 663) /w:[ 12 -1 11 18 ]
  //: joint g39 (w1) @(-76, 103) /w:[ 13 -1 14 16 ]
  myAND2 g195 (.A(w198), .B(w144), .Out(w201));   //: @(-747, 2090) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>0 Ti1>29 Bo0<1 ]
  //: joint g205 (w144) @(-330, 2029) /w:[ 8 -1 7 22 ]
  assign w154 = A[4]; //: TAP g179 @(-243,1666) /sn:0 /R:1 /w:[ 1 132 131 ] /ss:1
  assign w18 = A[6]; //: TAP g107 @(-207,623) /sn:0 /R:1 /w:[ 0 82 81 ] /ss:1
  FA g52 (.A(w11), .B(w24), .Cin(w27), .Cout(w33), .S(w34));   //: @(241, 518) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]
  myAND2 g231 (.B(w177), .A(w230), .Out(w234));   //: @(-872, 2471) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>29 Ti1>0 Bo0<1 ]
  FA g221 (.A(w200), .B(w196), .Cin(w222), .Cout(w227), .S(w228));   //: @(-671, 2237) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  assign w144 = B[6]; //: TAP g201 @(812,2029) /sn:0 /R:2 /w:[ 15 14 13 ] /ss:0
  assign w77 = A[4]; //: TAP g14 @(162,58) /sn:0 /R:1 /w:[ 1 55 56 ] /ss:1
  assign w12 = A[4]; //: TAP g44 @(91,299) /sn:0 /R:1 /w:[ 0 40 39 ] /ss:1
  myAND2 g47 (.A(w41), .B(w7), .Out(w8));   //: @(-269, 350) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<0 ]
  FA g247 (.A(w233), .B(w229), .Cin(w255), .Cout(w260), .S(w261));   //: @(-789, 2616) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g105 (w31) @(-308, 992) /w:[ 2 -1 1 28 ]
  FA g84 (.A(w58), .B(w57), .Cin(w60), .Cout(w61), .S(w63));   //: @(153, 894) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]
  //: joint g236 (w177) @(-180, 2434) /w:[ 12 -1 11 18 ]
  //: joint g23 (w1) @(124, 103) /w:[ 9 -1 10 20 ]
  FA g249 (.A(w237), .B(w239), .Cin(w265), .Cout(w270), .S(w271));   //: @(-1094, 2616) /sz:(90, 88) /sn:0 /p:[ Ti0>1 Ti1>0 Ri0>1 Lo0<1 Bo0<1 ]
  assign w81 = A[6]; //: TAP g116 @(-258,987) /sn:0 /R:1 /w:[ 1 100 99 ] /ss:1
  //: joint g40 (A) @(-284, 60) /w:[ 48 -1 66 47 ]
  myAND2 g93 (.B(w31), .A(w52), .Out(w70));   //: @(62, 1026) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>23 Ti1>0 Bo0<1 ]
  FA g54 (.A(w17), .B(w28), .Cin(w35), .Cout(w40), .S(w66));   //: @(19, 518) /sz:(90, 88) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  myAND2 g167 (.B(w136), .A(w169), .Out(w173));   //: @(-690, 1719) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<0 ]
  assign w92 = A[2]; //: TAP g46 @(312,299) /sn:0 /R:1 /w:[ 1 36 35 ] /ss:1
  //: IN g0 (A) @(-332,60) /sn:0 /w:[ 67 ]
  myAND2 g26 (.A(w94), .B(w7), .Out(w16));   //: @(376, 350) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>0 Ti1>19 Bo0<1 ]
  myAND2 g228 (.B(w177), .A(w215), .Out(w219));   //: @(-469, 2471) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>23 Ti1>0 Bo0<1 ]
  assign w165 = A[0]; //: TAP g224 @(-12,2392) /sn:0 /R:1 /w:[ 1 15 16 ] /ss:1
  assign w235 = A[7]; //: TAP g233 @(-975,2392) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  assign w111 = A[2]; //: TAP g136 @(121,1321) /sn:0 /R:1 /w:[ 1 110 109 ] /ss:1
  MyHA g173 (.B(w126), .A(w142), .cout(w149), .S(w155));   //: @(163, 1865) /sz:(107, 86) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<1 ]
  myAND2 g190 (.A(w170), .B(w144), .Out(w176));   //: @(-86, 2090) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>0 Ti1>19 Bo0<1 ]
  myAND2 g61 (.B(w4), .A(w97), .Out(w64));   //: @(78, 723) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>23 Ti1>0 Bo0<1 ]
  FA g220 (.A(w195), .B(w191), .Cin(w217), .Cout(w222), .S(w223));   //: @(-533, 2238) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  FA g86 (.A(w46), .B(w56), .Cin(w68), .Cout(w73), .S(w74));   //: @(-73, 895) /sz:(90, 88) /sn:0 /p:[ Ti0>1 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  //: joint g34 (w7) @(395, 268) /w:[ 12 -1 11 18 ]
  assign w3 = A[0]; //: TAP g3 @(646,59) /sn:0 /R:1 /w:[ 1 63 64 ] /ss:1
  assign w226 = {w221, w187, w155, w120, w103, w42, w22, w2}; //: CONCAT g250  @(-30,2970) /sn:0 /R:3 /w:[ 1 0 0 0 0 0 0 0 1 ] /dr:1 /tp:0 /drp:1
  myAND2 g65 (.B(w4), .A(w25), .Out(w65));   //: @(-371, 723) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Bo0<1 ]
  assign w100 = A[0]; //: TAP g110 @(424,972) /sn:0 /R:1 /w:[ 1 88 87 ] /ss:1
  myAND2 g59 (.B(w4), .A(w93), .Out(w43));   //: @(294, 723) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>19 Ti1>1 Bo0<1 ]
  //: joint g147 (w98) @(-140, 1353) /w:[ 6 -1 5 24 ]
  FA g156 (.A(w138), .B(w135), .Cin(w161), .Cout(w166), .S(w167));   //: @(-445, 1539) /sz:(90, 88) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]
  FA g153 (.A(w123), .B(w119), .Cin(w146), .Cout(w151), .S(w152));   //: @(-80, 1539) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  assign w31 = B[3]; //: TAP g98 @(812,992) /sn:0 /R:2 /w:[ 15 8 7 ] /ss:0
  myAND2 g96 (.B(w31), .A(w81), .Out(w85));   //: @(-327, 1026) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>29 Ti1>0 Bo0<1 ]
  assign w29 = A[2]; //: TAP g16 @(384,58) /sn:0 /R:1 /w:[ 1 59 60 ] /ss:1
  FA g183 (.A(w152), .B(w148), .Cin(w174), .Cout(w179), .S(w180));   //: @(-97, 1861) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  FA g122 (.A(w79), .B(w75), .Cin(w117), .Cout(w122), .S(w123));   //: @(-121, 1185) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  assign w93 = A[1]; //: TAP g78 @(350,623) /sn:0 /R:1 /w:[ 0 72 71 ] /ss:1
  FA g87 (.A(w51), .B(w59), .Cin(w73), .Cout(w78), .S(w79));   //: @(-186, 895) /sz:(90, 88) /sn:0 /p:[ Ti0>1 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  //: joint g171 (w136) @(88, 1686) /w:[ 12 -1 11 18 ]
  myAND2 g129 (.A(w116), .B(w98), .Out(w119));   //: @(-42, 1375) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>0 Ti1>23 Bo0<1 ]
  assign w225 = A[5]; //: TAP g258 @(-673,2392) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  FA g244 (.A(w218), .B(w214), .Cin(w240), .Cout(w245), .S(w246));   //: @(-385, 2616) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  //: joint g143 (w98) @(319, 1353) /w:[ 14 -1 13 16 ]
  //: joint g69 (w4) @(204, 663) /w:[ 10 -1 9 20 ]
  FA g245 (.A(w223), .B(w219), .Cin(w245), .Cout(w250), .S(w251));   //: @(-513, 2616) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<1 ]
  FA g119 (.A(w63), .B(w44), .Cin(w102), .Cout(w107), .S(w108));   //: @(246, 1185) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  assign w82 = A[3]; //: TAP g15 @(273,58) /sn:0 /R:1 /w:[ 1 57 58 ] /ss:1
  myAND2 g162 (.B(w136), .A(w110), .Out(w148));   //: @(-60, 1719) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>21 Ti1>1 Bo0<1 ]
  myAND2 g127 (.A(w106), .B(w98), .Out(w109));   //: @(175, 1374) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>0 Ti1>19 Bo0<0 ]
  //: joint g67 (w4) @(441, 663) /w:[ 14 -1 13 16 ]
  myAND2 g131 (.A(w129), .B(w98), .Out(w130));   //: @(-283, 1380) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>0 Ti1>27 Bo0<1 ]
  assign w48 = A[5]; //: TAP g43 @(-7,299) /sn:0 /R:1 /w:[ 0 42 41 ] /ss:1
  myAND2 g62 (.B(w4), .A(w72), .Out(w56));   //: @(-26, 723) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>25 Ti1>1 Bo0<1 ]
  FA g88 (.A(w55), .B(w62), .Cin(w78), .Cout(w83), .S(w125));   //: @(-310, 895) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<1 ]
  //: joint g104 (w31) @(-181, 992) /w:[ 4 -1 3 26 ]
  FA g188 (.A(w171), .B(w173), .Cin(w199), .Cout(w204), .S(w205));   //: @(-738, 1857) /sz:(90, 88) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]
  myAND2 g63 (.B(w4), .A(w15), .Out(w59));   //: @(-145, 723) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>27 Ti1>1 Bo0<1 ]
  assign w121 = A[4]; //: TAP g138 @(-102,1321) /sn:0 /R:1 /w:[ 1 114 113 ] /ss:1
  assign w220 = A[4]; //: TAP g257 @(-538,2392) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  //: joint g109 (A) @(656, 980) /w:[ -1 24 86 23 ]
  //: joint g175 (w136) @(-418, 1686) /w:[ 4 -1 3 26 ]
  assign w177 = B[7]; //: TAP g234 @(812,2434) /sn:0 /R:2 /w:[ 15 16 15 ] /ss:0
  myAND2 g133 (.A(w139), .B(w98), .Out(w140));   //: @(-526, 1378) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<0 ]
  FA g56 (.A(w23), .B(w32), .Cin(w45), .Cout(w50), .S(w51));   //: @(-216, 519) /sz:(90, 88) /sn:0 /p:[ Ti0>1 Ti1>0 Ri0>1 Lo0<0 Bo0<0 ]
  myAND2 g5 (.B(w1), .A(w29), .Out(w19));   //: @(328, 128) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>25 Ti1>0 Bo0<0 ]
  myAND2 g95 (.B(w31), .A(w76), .Out(w80));   //: @(-200, 1026) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>27 Ti1>0 Bo0<1 ]
  myAND2 g92 (.B(w31), .A(w87), .Out(w49));   //: @(171, 1026) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>21 Ti1>1 Bo0<0 ]
  //: joint g24 (w1) @(21, 103) /w:[ 11 -1 12 18 ]
  FA g85 (.A(w66), .B(w64), .Cin(w61), .Cout(w68), .S(w69));   //: @(32, 895) /sz:(90, 88) /sn:0 /p:[ Ti0>1 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  assign w198 = A[6]; //: TAP g214 @(-689,1994) /sn:0 /R:1 /w:[ 1 154 153 ] /ss:1
  assign w178 = A[2]; //: TAP g210 @(-161,1995) /sn:0 /R:1 /w:[ 1 146 145 ] /ss:1
  //: joint g101 (w31) @(190, 992) /w:[ 10 -1 9 20 ]
  myAND2 g60 (.B(w4), .A(w91), .Out(w57));   //: @(185, 723) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>21 Ti1>0 Bo0<0 ]
  assign w253 = {w270, w271, w266, w261, w256, w251, w246, w241}; //: CONCAT g251  @(-261,2970) /sn:0 /R:3 /w:[ 1 0 0 0 1 0 0 0 0 ] /dr:1 /tp:0 /drp:1
  //: joint g204 (w144) @(-199, 2029) /w:[ 10 -1 9 20 ]
  FA g185 (.A(w162), .B(w158), .Cin(w181), .Cout(w189), .S(w190));   //: @(-338, 1858) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  //: joint g35 (w7) @(274, 268) /w:[ 10 -1 9 20 ]
  myAND2 g126 (.A(w101), .B(w98), .Out(w104));   //: @(301, 1373) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>0 Ti1>17 Bo0<0 ]
  //: joint g170 (w136) @(215, 1686) /w:[ 14 -1 13 16 ]
  FA g120 (.A(w69), .B(w49), .Cin(w107), .Cout(w112), .S(w113));   //: @(140, 1185) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g235 (w177) @(-50, 2434) /w:[ 14 -1 13 16 ]
  assign w4 = B[2]; //: TAP g66 @(812,663) /sn:0 /R:2 /w:[ 15 6 5 ] /ss:0
  myAND2 g97 (.B(w31), .A(w86), .Out(w90));   //: @(-448, 1026) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<1 ]
  FA g184 (.A(w157), .B(w153), .Cin(w179), .Cout(w181), .S(w185));   //: @(-227, 1859) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  //: joint g260 (A) @(656, 1995) /w:[ -1 18 140 17 ]
  myAND2 g226 (.B(w177), .A(w197), .Out(w209));   //: @(-199, 2471) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>19 Ti1>0 Bo0<1 ]
  assign w47 = A[6]; //: TAP g12 @(-39,58) /sn:0 /R:1 /w:[ 1 51 52 ] /ss:1
  assign w1 = B[0]; //: TAP g18 @(812,103) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:0
  //: joint g239 (w177) @(-575, 2434) /w:[ 6 -1 5 24 ]
  //: joint g108 (A) @(657, 625) /w:[ -1 26 68 25 ]
  myAND2 g191 (.A(w178), .B(w144), .Out(w182));   //: @(-218, 2090) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>0 Ti1>21 Bo0<1 ]
  FA g219 (.A(w190), .B(w186), .Cin(w212), .Cout(w217), .S(w218));   //: @(-405, 2238) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  MyHA g242 (.B(w192), .A(w208), .cout(w216), .S(w221));   //: @(-115, 2606) /sz:(107, 86) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<1 ]
  assign w101 = A[0]; //: TAP g134 @(359,1321) /sn:0 /R:1 /w:[ 1 106 105 ] /ss:1
  myAND2 g4 (.B(w1), .A(w6), .Out(w13));   //: @(462, 128) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>27 Ti1>0 Bo0<0 ]
  FA g154 (.A(w128), .B(w124), .Cin(w151), .Cout(w156), .S(w157));   //: @(-200, 1539) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  //: joint g237 (w177) @(-314, 2434) /w:[ 10 -1 9 20 ]
  myAND2 g58 (.B(w4), .A(w95), .Out(w0));   //: @(422, 723) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>17 Ti1>1 Bo0<0 ]
  FA g186 (.A(w167), .B(w163), .Cin(w189), .Cout(w194), .S(w195));   //: @(-481, 1855) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  assign w87 = A[2]; //: TAP g112 @(228,978) /sn:0 /R:1 /w:[ 0 92 91 ] /ss:1
  assign w25 = A[7]; //: TAP g76 @(-314,623) /sn:0 /R:1 /w:[ 0 84 83 ] /ss:1
  assign w184 = A[3]; //: TAP g211 @(-293,1995) /sn:0 /R:1 /w:[ 1 148 147 ] /ss:1
  FA g157 (.A(w137), .B(w140), .Cin(w166), .Cout(w171), .S(w172));   //: @(-564, 1538) /sz:(90, 88) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]
  myAND2 g163 (.B(w136), .A(w150), .Out(w153));   //: @(-184, 1719) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>23 Ti1>0 Bo0<1 ]
  //: joint g238 (w177) @(-450, 2434) /w:[ 8 -1 7 22 ]
  assign w230 = A[6]; //: TAP g259 @(-815,2392) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  myAND2 g64 (.B(w4), .A(w18), .Out(w62));   //: @(-264, 718) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>29 Ti1>1 Bo0<1 ]
  myAND2 g166 (.B(w136), .A(w164), .Out(w168));   //: @(-568, 1719) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>29 Ti1>0 Bo0<1 ]
  FA g121 (.A(w74), .B(w70), .Cin(w112), .Cout(w117), .S(w118));   //: @(12, 1185) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g206 (w144) @(-462, 2029) /w:[ 6 -1 5 24 ]
  //: joint g241 (w177) @(-853, 2434) /w:[ 2 -1 1 28 ]
  myAND2 g28 (.B(w7), .A(w9), .Out(w26));   //: @(139, 350) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>23 Ti1>1 Bo0<1 ]
  myAND2 g225 (.B(w177), .A(w165), .Out(w192));   //: @(-69, 2471) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>17 Ti1>0 Bo0<0 ]
  myAND2 g6 (.B(w1), .A(w82), .Out(w11));   //: @(216, 128) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>23 Ti1>0 Bo0<1 ]
  assign w159 = A[5]; //: TAP g177 @(-380,1666) /sn:0 /R:1 /w:[ 1 134 133 ] /ss:1
  myAND2 g192 (.A(w184), .B(w144), .Out(w186));   //: @(-348, 2090) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>0 Ti1>23 Bo0<1 ]
  //: joint g208 (w144) @(-728, 2029) /w:[ 2 -1 1 28 ]
  myAND2 g7 (.B(w1), .A(w77), .Out(w14));   //: @(105, 128) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>21 Ti1>0 Bo0<0 ]
  FA g53 (.A(w14), .B(w26), .Cin(w33), .Cout(w35), .S(w58));   //: @(122, 518) /sz:(90, 88) /sn:0 /p:[ Ti0>1 Ti1>0 Ri0>0 Lo0<0 Bo0<1 ]
  //: joint g149 (w98) @(-382, 1353) /w:[ 2 -1 1 28 ]
  //: joint g207 (w144) @(-589, 2029) /w:[ 4 -1 3 26 ]
  //: joint g48 (w7) @(-148, 268) /w:[ 2 -1 1 28 ]
  assign w110 = A[2]; //: TAP g200 @(-3,1666) /sn:0 /R:1 /w:[ 0 128 127 ] /ss:1
  myAND2 g25 (.A(w96), .B(w7), .Out(w10));   //: @(512, 350) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>0 Ti1>17 Bo0<0 ]
  assign w6 = A[1]; //: TAP g17 @(520,58) /sn:0 /R:1 /w:[ 1 61 62 ] /ss:1
  myAND2 g29 (.B(w7), .A(w12), .Out(w28));   //: @(35, 350) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>25 Ti1>1 Bo0<0 ]
  assign w15 = A[5]; //: TAP g106 @(-88,623) /sn:0 /R:1 /w:[ 0 80 79 ] /ss:1
  FA g83 (.A(w34), .B(w43), .Cin(w38), .Cout(w60), .S(w53));   //: @(263, 895) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<0 Bo0<0 ]
  //: joint g174 (w136) @(-281, 1686) /w:[ 6 -1 5 24 ]
  //: joint g100 (w31) @(298, 992) /w:[ 12 -1 11 18 ]
  myAND2 g94 (.B(w31), .A(w71), .Out(w75));   //: @(-70, 1026) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>25 Ti1>0 Bo0<1 ]
  assign w97 = A[3]; //: TAP g80 @(134,623) /sn:0 /R:1 /w:[ 1 76 75 ] /ss:1
  myAND2 g193 (.A(w188), .B(w144), .Out(w191));   //: @(-481, 2090) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>0 Ti1>25 Bo0<1 ]
  //: joint g202 (w144) @(65, 2029) /w:[ 14 -1 13 16 ]
  FA g248 (.A(w238), .B(w234), .Cin(w260), .Cout(w265), .S(w266));   //: @(-952, 2616) /sz:(90, 88) /sn:0 /p:[ Ti0>1 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  //: OUT g253 (Out) @(-148,3092) /sn:0 /R:3 /w:[ 1 ]
  //: joint g21 (w1) @(347, 103) /w:[ 5 -1 6 24 ]
  //: joint g159 (A) @(656, 1666) /w:[ -1 20 122 19 ]
  //: joint g172 (w136) @(-41, 1686) /w:[ 10 -1 9 20 ]
  myAND2 g232 (.B(w177), .A(w235), .Out(w239));   //: @(-1031, 2471) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<1 ]
  assign w41 = A[7]; //: TAP g41 @(-212,299) /sn:0 /R:1 /w:[ 1 46 45 ] /ss:1
  assign w139 = A[6]; //: TAP g141 @(-468,1321) /sn:0 /R:1 /w:[ 1 120 119 ] /ss:1
  FA g155 (.A(w133), .B(w130), .Cin(w156), .Cout(w161), .S(w162));   //: @(-328, 1540) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  assign w215 = A[3]; //: TAP g256 @(-412,2392) /sn:0 /R:1 /w:[ 1 9 10 ] /ss:1
  FA g123 (.A(w125), .B(w80), .Cin(w122), .Cout(w127), .S(w128));   //: @(-249, 1185) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  FA g151 (.A(w113), .B(w109), .Cin(w115), .Cout(w141), .S(w142));   //: @(155, 1543) /sz:(90, 88) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<0 ]
  myAND2 g90 (.B(w31), .A(w100), .Out(w36));   //: @(377, 1026) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>17 Ti1>0 Bo0<0 ]
  FA g222 (.A(w205), .B(w201), .Cin(w227), .Cout(w232), .S(w233));   //: @(-806, 2237) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  MyHA g82 (.B(w0), .A(w37), .cout(w38), .S(w42));   //: @(425, 877) /sz:(107, 86) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<1 ]
  myAND2 g128 (.A(w111), .B(w98), .Out(w114));   //: @(65, 1374) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>0 Ti1>21 Bo0<1 ]
  FA g243 (.A(w213), .B(w209), .Cin(w216), .Cout(w240), .S(w241));   //: @(-251, 2616) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<0 Bo0<1 ]
  //: joint g33 (w7) @(531, 268) /w:[ 14 -1 13 16 ]
  myAND2 g91 (.B(w31), .A(w99), .Out(w44));   //: @(279, 1026) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>19 Ti1>0 Bo0<1 ]
  assign w94 = A[1]; //: TAP g49 @(432,298) /sn:0 /R:1 /w:[ 1 34 33 ] /ss:1
  assign w116 = A[3]; //: TAP g137 @(13,1321) /sn:0 /R:1 /w:[ 1 112 111 ] /ss:1
  assign w105 = A[0]; //: TAP g198 @(254,1666) /sn:0 /R:1 /w:[ 1 124 123 ] /ss:1
  FA g51 (.A(w19), .B(w16), .Cin(w5), .Cout(w27), .S(w37));   //: @(363, 518) /sz:(90, 88) /sn:0 /p:[ Ti0>1 Ti1>0 Ri0>0 Lo0<0 Bo0<0 ]
  //: joint g158 (A) @(656, 1323) /w:[ -1 22 104 21 ]
  FA g89 (.A(w54), .B(w65), .Cin(w83), .Cout(w88), .S(w89));   //: @(-428, 895) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<0 Bo0<1 ]
  FA g217 (.A(w180), .B(w176), .Cin(w183), .Cout(w207), .S(w208));   //: @(-141, 2238) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<0 ]
  assign w95 = A[0]; //: TAP g77 @(479,623) /sn:0 /R:1 /w:[ 0 70 69 ] /ss:1
  myAND2 g2 (.B(w1), .A(w3), .Out(w2));   //: @(590, 128) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>29 Ti1>0 Bo0<0 ]
  assign w193 = A[5]; //: TAP g213 @(-551,1994) /sn:0 /R:1 /w:[ 1 152 151 ] /ss:1
  //: joint g148 (w98) @(-264, 1353) /w:[ 4 -1 3 26 ]
  assign Out = {w253, w226}; //: CONCAT g252  @(-148,3050) /sn:0 /R:3 /w:[ 0 0 0 ] /dr:1 /tp:0 /drp:1
  //: joint g203 (w144) @(-67, 2029) /w:[ 12 -1 11 18 ]
  //: joint g72 (w4) @(-114, 663) /w:[ 4 -1 3 26 ]
  //: joint g99 (w31) @(395, 992) /w:[ 14 -1 13 16 ]
  myAND2 g161 (.B(w136), .A(w131), .Out(w143));   //: @(69, 1719) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>19 Ti1>0 Bo0<1 ]
  FA g182 (.A(w147), .B(w143), .Cin(w149), .Cout(w174), .S(w175));   //: @(34, 1864) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<0 Bo0<0 ]
  myAND2 g196 (.A(w203), .B(w144), .Out(w206));   //: @(-878, 2090) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<1 ]
  //: joint g103 (w31) @(-51, 992) /w:[ 6 -1 5 24 ]
  FA g152 (.A(w118), .B(w114), .Cin(w141), .Cout(w146), .S(w147));   //: @(37, 1541) /sz:(90, 88) /sn:0 /p:[ Ti0>1 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  myAND2 g189 (.A(w145), .B(w144), .Out(w160));   //: @(46, 2090) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>0 Ti1>17 Bo0<0 ]
  FA g246 (.A(w228), .B(w224), .Cin(w250), .Cout(w255), .S(w256));   //: @(-651, 2616) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<0 Bo0<1 ]
  assign w210 = A[2]; //: TAP g255 @(-276,2392) /sn:0 /R:1 /w:[ 1 11 12 ] /ss:1
  myAND2 g10 (.B(w1), .A(w21), .Out(w23));   //: @(-201, 128) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>15 Ti1>0 Bo0<0 ]
  assign w188 = A[4]; //: TAP g212 @(-424,1995) /sn:0 /R:1 /w:[ 1 150 149 ] /ss:1
  myAND2 g27 (.B(w7), .A(w92), .Out(w24));   //: @(255, 350) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>21 Ti1>0 Bo0<0 ]
  assign w7 = B[1]; //: TAP g32 @(812,268) /sn:0 /R:2 /w:[ 15 4 3 ] /ss:0
  assign w131 = A[1]; //: TAP g199 @(126,1666) /sn:0 /R:1 /w:[ 1 126 125 ] /ss:1
  //: joint g102 (w31) @(81, 992) /w:[ 8 -1 7 22 ]
  FA g187 (.A(w172), .B(w168), .Cin(w194), .Cout(w199), .S(w200));   //: @(-607, 1858) /sz:(90, 88) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  //: joint g240 (w177) @(-709, 2434) /w:[ 4 -1 3 26 ]
  MyHA g57 (.B(w50), .A(w8), .cout(w54), .S(w55));   //: @(-354, 505) /sz:(107, 86) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<1 ]
  myAND2 g9 (.B(w1), .A(w47), .Out(w20));   //: @(-95, 128) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>17 Ti1>0 Bo0<1 ]
  //: joint g71 (w4) @(-7, 663) /w:[ 6 -1 5 24 ]
  assign w98 = B[4]; //: TAP g142 @(812,1353) /sn:0 /R:2 /w:[ 15 10 9 ] /ss:0
  //: joint g145 (w98) @(84, 1353) /w:[ 10 -1 9 20 ]
  //: joint g73 (w4) @(-216, 663) /w:[ 2 -1 1 28 ]
  assign w39 = A[6]; //: TAP g42 @(-110,299) /sn:0 /R:1 /w:[ 0 44 43 ] /ss:1
  assign w150 = A[3]; //: TAP g180 @(-128,1666) /sn:0 /R:1 /w:[ 1 130 129 ] /ss:1
  assign w96 = A[0]; //: TAP g74 @(569,299) /sn:0 /R:1 /w:[ 1 32 31 ] /ss:1
  //: joint g181 (w136) @(-169, 1686) /w:[ 8 -1 7 22 ]
  assign w169 = A[7]; //: TAP g168 @(-633,1666) /sn:0 /R:1 /w:[ 1 138 137 ] /ss:1
  assign w91 = A[2]; //: TAP g79 @(240,623) /sn:0 /R:1 /w:[ 1 74 73 ] /ss:1
  assign w86 = A[7]; //: TAP g117 @(-403,978) /sn:0 /R:1 /w:[ 1 102 101 ] /ss:1
  myAND2 g194 (.A(w193), .B(w144), .Out(w196));   //: @(-608, 2090) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>0 Ti1>27 Bo0<1 ]
  assign w203 = A[7]; //: TAP g215 @(-821,1994) /sn:0 /R:1 /w:[ 1 156 155 ] /ss:1
  MyHA g216 (.B(w160), .A(w175), .cout(w183), .S(w187));   //: @(13, 2230) /sz:(107, 86) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<0 Bo0<1 ]
  //: joint g36 (w7) @(158, 268) /w:[ 8 -1 7 22 ]
  FA g125 (.A(w88), .B(w90), .Cin(w132), .Cout(w137), .S(w138));   //: @(-494, 1185) /sz:(90, 88) /sn:0 /p:[ Ti0>1 Ti1>0 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g144 (w98) @(194, 1353) /w:[ 12 -1 11 18 ]
  assign w164 = A[6]; //: TAP g178 @(-513,1666) /sn:0 /R:1 /w:[ 1 136 135 ] /ss:1
  assign w72 = A[4]; //: TAP g81 @(30,623) /sn:0 /R:1 /w:[ 0 78 77 ] /ss:1
  //: joint g22 (w1) @(235, 103) /w:[ 7 -1 8 22 ]
  //: joint g70 (w4) @(97, 663) /w:[ 8 -1 7 22 ]
  assign w9 = A[3]; //: TAP g45 @(196,299) /sn:0 /R:1 /w:[ 0 38 37 ] /ss:1
  assign w170 = A[1]; //: TAP g209 @(-29,1993) /sn:0 /R:1 /w:[ 1 144 143 ] /ss:1
  assign w71 = A[4]; //: TAP g114 @(-14,978) /sn:0 /R:1 /w:[ 1 96 95 ] /ss:1
  myAND2 g229 (.B(w177), .A(w220), .Out(w224));   //: @(-594, 2471) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>25 Ti1>0 Bo0<1 ]
  myAND2 g30 (.B(w7), .A(w48), .Out(w30));   //: @(-64, 350) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>27 Ti1>1 Bo0<1 ]
  myAND2 g164 (.B(w136), .A(w154), .Out(w158));   //: @(-300, 1719) /sz:(79, 103) /R:3 /sn:0 /p:[ Ti0>25 Ti1>0 Bo0<1 ]
  MyHA g118 (.B(w36), .A(w53), .cout(w102), .S(w103));   //: @(369, 1179) /sz:(107, 86) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<0 Bo0<1 ]

endmodule
//: /netlistEnd

//: /netlistBegin FlipFlopDLS
module FlipFlopDLS(Clk, D, Y);
//: interface  /sz:(116, 96) /bd:[ Li0>D(24/96) Bi0>Clk(62/116) Ro0<Y(21/96) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input Clk;    //: /sn:0 {0}(388,329)(399,329)(399,268){1}
input D;    //: /sn:0 {0}(125,187)(176,187){1}
//: {2}(180,187)(309,187)(309,207)(355,207){3}
//: {4}(178,189)(178,245)(186,245){5}
output Y;    //: /sn:0 {0}(443,208)(534,208)(534,206)(549,206){1}
wire w1;    //: /sn:0 {0}(355,254)(303,254)(303,263)(238,263){1}
//: enddecls

  //: IN g4 (Clk) @(386,329) /sn:0 /w:[ 0 ]
  //: joint g3 (D) @(178, 187) /w:[ 2 -1 1 4 ]
  //: IN g2 (D) @(123,187) /sn:0 /w:[ 0 ]
  myINV g1 (.In(D), .Out(w1));   //: @(187, 233) /sz:(50, 46) /sn:0 /p:[ Li0>5 Ro0<1 ]
  //: OUT g5 (Y) @(546,206) /sn:0 /w:[ 1 ]
  FlipFlopSR g0 (.R(w1), .S(D), .Clk(Clk), .Y(Y));   //: @(356, 192) /sz:(86, 75) /sn:0 /p:[ Li0>0 Li1>3 Bi0>1 Ro0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin FlipFlopSR
module FlipFlopSR(R, S, Y, Clk);
//: interface  /sz:(86, 75) /bd:[ Li0>S(15/75) Li1>R(62/75) Bi0>Clk(43/86) Ro0<Y(16/75) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input R;    //: /sn:0 {0}(95,259)(188,259)(188,281)(218,281){1}
input Clk;    //: /sn:0 {0}(218,243)(166,243)(166,235)(156,235){1}
//: {2}(154,233)(154,174)(203,174){3}
//: {4}(154,237)(154,362)(168,362)(168,375)(158,375){5}
input S;    //: /sn:0 {0}(116,127)(173,127)(173,136)(203,136){1}
output Y;    //: /sn:0 {0}(607,220)(524,220)(524,219)(509,219){1}
wire w3;    //: /sn:0 {0}(524,165)(509,165){1}
wire w0;    //: /sn:0 {0}(406,163)(359,163)(359,155)(308,155){1}
wire w1;    //: /sn:0 {0}(406,218)(396,218)(396,262)(323,262){1}
//: enddecls

  //: IN g4 (R) @(93,259) /sn:0 /w:[ 0 ]
  //: IN g3 (S) @(114,127) /sn:0 /w:[ 0 ]
  myAND2 g2 (.B(R), .A(Clk), .Out(w1));   //: @(219, 222) /sz:(103, 79) /sn:0 /p:[ Li0>1 Li1>0 Ro0<1 ]
  myAND2 g1 (.B(Clk), .A(S), .Out(w0));   //: @(204, 115) /sz:(103, 79) /sn:0 /p:[ Li0>3 Li1>1 Ro0<1 ]
  //: joint g6 (Clk) @(154, 235) /w:[ 1 2 -1 4 ]
  //: OUT g7 (Y) @(604,220) /sn:0 /w:[ 0 ]
  //: IN g5 (Clk) @(156,375) /sn:0 /w:[ 5 ]
  latchSR g0 (.R(w1), .S(w0), .Y(Y), .Y1(w3));   //: @(407, 138) /sz:(101, 105) /sn:0 /p:[ Li0>0 Li1>0 Ri0>1 Ro0<1 ]

endmodule
//: /netlistEnd

//: /netlistBegin MyHA
module MyHA(cout, B, A, S);
//: interface  /sz:(107, 86) /bd:[ Ti0>A(89/107) Ti1>B(28/107) Lo0<cout(41/86) Bo0<S(54/107) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input B;    //: /sn:0 {0}(471,382)(277,382)(277,142){1}
//: {2}(279,140)(376,140)(376,135)(426,135){3}
//: {4}(275,140)(213,140)(213,296)(103,296){5}
input A;    //: /sn:0 {0}(471,344)(376,344)(376,118){1}
//: {2}(378,116)(405,116)(405,115)(426,115){3}
//: {4}(374,116)(152,116)(152,179)(116,179){5}
output S;    //: /sn:0 {0}(808,122)(615,122)(615,129)(515,129){1}
output cout;    //: /sn:0 {0}(576,363)(651,363)(651,354)(848,354){1}
//: enddecls

  //: OUT g4 (cout) @(845,354) /sn:0 /w:[ 1 ]
  myEXOR g8 (.A(A), .B(B), .Out(S));   //: @(427, 99) /sz:(87, 60) /sn:0 /p:[ Li0>3 Li1>3 Ro0<1 ]
  //: IN g3 (B) @(101,296) /sn:0 /w:[ 5 ]
  //: IN g2 (A) @(114,179) /sn:0 /w:[ 5 ]
  //: joint g1 (A) @(376, 116) /w:[ 2 -1 4 1 ]
  //: joint g6 (B) @(277, 140) /w:[ 2 -1 4 1 ]
  //: OUT g5 (S) @(805,122) /sn:0 /w:[ 0 ]
  myAND2 g0 (.B(B), .A(A), .Out(cout));   //: @(472, 323) /sz:(103, 79) /sn:0 /p:[ Li0>0 Li1>0 Ro0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin MYADDER18
module MYADDER18(A, Cout, Cin, S, B);
//: interface  /sz:(164, 142) /bd:[ Ti0>B[17:0](116/164) Ti1>A[17:0](23/164) Ri0>Cin(59/142) Lo0<Cout(62/142) Bo0<S[17:0](68/164) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [17:0] B;    //: /sn:0 {0}(#:1330,103)(1204,103){1}
//: {2}(1203,103)(1003,103){3}
//: {4}(1002,103)(793,103){5}
//: {6}(792,103)(653,103){7}
//: {8}(652,103)(291,103){9}
//: {10}(290,103)(#:48,103){11}
input [17:0] A;    //: /sn:0 {0}(#:1336,66)(1145,66){1}
//: {2}(1144,66)(944,66){3}
//: {4}(943,66)(736,66){5}
//: {6}(735,66)(594,66){7}
//: {8}(593,66)(223,66){9}
//: {10}(222,66)(#:54,66){11}
output Cout;    //: /sn:0 {0}(185,227)(99,227)(99,240)(89,240){1}
input Cin;    //: /sn:0 {0}(1330,257)(1271,257)(1271,244)(1253,244){1}
output [17:0] S;    //: /sn:0 {0}(#:1229,404)(1362,404){1}
wire [3:0] w6;    //: /sn:0 {0}(653,107)(#:653,117)(539,117)(539,223){1}
wire [3:0] w7;    //: /sn:0 {0}(#:723,229)(723,82)(736,82)(736,70){1}
wire [1:0] w16;    //: /sn:0 {0}(291,107)(#:291,137)(276,137)(276,207){1}
wire [3:0] w14;    //: /sn:0 {0}(#:513,265)(513,394)(#:1223,394){1}
wire [3:0] w15;    //: /sn:0 {0}(#:977,269)(977,414)(1223,414){1}
wire w4;    //: /sn:0 {0}(588,236)(665,236)(665,242)(686,242){1}
wire [3:0] w0;    //: /sn:0 {0}(#:1145,70)(1145,187)(1143,187)(1143,231){1}
wire [3:0] w3;    //: /sn:0 {0}(1178,273)(1178,424)(#:1223,424){1}
wire w21;    //: /sn:0 {0}(1106,244)(1060,244)(1060,240)(1052,240){1}
wire [1:0] w23;    //: /sn:0 {0}(251,261)(251,384)(#:1223,384){1}
wire [3:0] w1;    //: /sn:0 {0}(#:1204,107)(1204,231){1}
wire [3:0] w8;    //: /sn:0 {0}(#:1003,227)(1003,107){1}
wire w18;    //: /sn:0 {0}(325,226)(431,226)(431,236)(441,236){1}
wire w22;    //: /sn:0 {0}(905,240)(843,240)(843,242)(833,242){1}
wire [1:0] w11;    //: /sn:0 {0}(#:223,70)(223,192)(219,192)(219,207){1}
wire [3:0] w2;    //: /sn:0 {0}(#:784,229)(784,119)(793,119)(793,107){1}
wire [3:0] w10;    //: /sn:0 {0}(#:758,271)(758,404)(#:1223,404){1}
wire [3:0] w13;    //: /sn:0 {0}(#:942,227)(942,78)(944,78)(944,70){1}
wire [3:0] w5;    //: /sn:0 {0}(594,70)(#:594,80)(478,80)(478,223){1}
//: enddecls

  //: IN g4 (A) @(52,66) /sn:0 /w:[ 11 ]
  assign w16 = B[17:16]; //: TAP g8 @(291,101) /sn:0 /R:1 /w:[ 0 10 9 ] /ss:1
  MYADDER4 g13 (.A(w13), .B(w8), .Cin(w21), .Cout(w22), .S(w15));   //: @(906, 228) /sz:(145, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<0 ]
  //: OUT g3 (Cout) @(92,240) /sn:0 /R:2 /w:[ 1 ]
  //: IN g2 (Cin) @(1332,257) /sn:0 /R:2 /w:[ 0 ]
  MYADDER4 g1 (.A(w5), .B(w6), .Cin(w4), .Cout(w18), .S(w14));   //: @(442, 224) /sz:(145, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]
  assign w2 = B[11:8]; //: TAP g16 @(793,101) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  //: OUT g11 (S) @(1359,404) /sn:0 /w:[ 1 ]
  assign S = {w23, w14, w10, w15, w3}; //: CONCAT g10  @(1228,404) /sn:0 /w:[ 0 1 1 1 1 1 ] /dr:0 /tp:0 /drp:1
  assign w0 = A[3:0]; //: TAP g19 @(1145,64) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  assign w11 = A[17:16]; //: TAP g6 @(223,64) /sn:0 /R:1 /w:[ 0 10 9 ] /ss:1
  assign w5 = A[15:12]; //: TAP g7 @(594,64) /sn:0 /R:1 /w:[ 0 8 7 ] /ss:1
  assign w6 = B[15:12]; //: TAP g9 @(653,101) /sn:0 /R:1 /w:[ 0 8 7 ] /ss:1
  assign w1 = B[3:0]; //: TAP g20 @(1204,101) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  assign w7 = A[11:8]; //: TAP g15 @(736,64) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  assign w13 = A[7:4]; //: TAP g17 @(944,64) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  MYADDER2 g14 (.A(w11), .B(w16), .Cin(w18), .Cout(Cout), .S(w23));   //: @(186, 208) /sz:(138, 52) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<0 Bo0<0 ]
  //: IN g5 (B) @(46,103) /sn:0 /w:[ 11 ]
  MYADDER4 g0 (.A(w0), .B(w1), .Cin(Cin), .Cout(w21), .S(w3));   //: @(1107, 232) /sz:(145, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  assign w8 = B[7:4]; //: TAP g18 @(1003,101) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  MYADDER4 g12 (.A(w7), .B(w2), .Cin(w22), .Cout(w4), .S(w10));   //: @(687, 230) /sz:(145, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin myAND2
module myAND2(Out, B, A);
//: interface  /sz:(103, 79) /bd:[ Li0>A(21/79) Li1>B(59/79) Ro0<Out(40/79) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input B;    //: /sn:0 {0}(212,195)(257,195){1}
input A;    //: /sn:0 {0}(257,167)(209,167){1}
output Out;    //: /sn:0 {0}(578,181)(505,181)(505,189)(480,189){1}
wire w2;    //: /sn:0 {0}(425,182)(422,182){1}
//: {2}(420,180)(420,171)(428,171){3}
//: {4}(418,182)(378,182){5}
//: enddecls

  //: OUT g4 (Out) @(575,181) /sn:0 /w:[ 0 ]
  myINV g3 (.In(w2), .Out(Out));   //: @(429, 159) /sz:(50, 46) /sn:0 /p:[ Li0>3 Ro0<1 ]
  myNAND2 g2 (.B(B), .A(A), .Out(w2));   //: @(258, 150) /sz:(119, 61) /sn:0 /p:[ Li0>1 Li1>0 Ro0<5 ]
  //: IN g1 (B) @(210,195) /sn:0 /w:[ 0 ]
  //: joint g5 (w2) @(420, 182) /w:[ 1 2 4 -1 ]
  //: IN g0 (A) @(207,167) /sn:0 /w:[ 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin MyCOMPLEMENT2
module MyCOMPLEMENT2(In, Out, minus, Cout);
//: interface  /sz:(138, 79) /bd:[ Li0>minus(63/79) Li1>In[17:0](36/79) To0<Cout(62/138) Ro0<Out[17:0](34/79) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [17:0] In;    //: /sn:0 {0}(#:2558,34)(2510,34){1}
//: {2}(2509,34)(2370,34){3}
//: {4}(2369,34)(2254,34){5}
//: {6}(2253,34)(2111,34){7}
//: {8}(2110,34)(1996,34){9}
//: {10}(1995,34)(1863,34){11}
//: {12}(1862,34)(1715,34){13}
//: {14}(1714,34)(1599,34){15}
//: {16}(1598,34)(1455,34){17}
//: {18}(1454,34)(1345,34){19}
//: {20}(1344,34)(1155,34){21}
//: {22}(1154,34)(1037,34){23}
//: {24}(1036,34)(917,34){25}
//: {26}(916,34)(785,34){27}
//: {28}(784,34)(668,34){29}
//: {30}(667,34)(544,34){31}
//: {32}(543,34)(334,34){33}
//: {34}(333,34)(105,34){35}
//: {36}(104,34)(#:46,34){37}
input minus;    //: /sn:0 {0}(2575,304)(2575,107)(2576,107)(2576,97){1}
//: {2}(2578,95)(2591,95)(2591,30){3}
//: {4}(2574,95)(2538,95){5}
//: {6}(2534,95)(2399,95){7}
//: {8}(2395,95)(2272,95){9}
//: {10}(2268,95)(2133,95){11}
//: {12}(2129,95)(2018,95){13}
//: {14}(2014,95)(1883,95){15}
//: {16}(1879,95)(1735,95){17}
//: {18}(1731,95)(1623,95){19}
//: {20}(1619,95)(1479,95){21}
//: {22}(1475,95)(1367,95){23}
//: {24}(1363,95)(1190,95){25}
//: {26}(1188,93)(1188,90)(1203,90)(1203,108){27}
//: {28}(1186,95)(1068,95){29}
//: {30}(1066,93)(1066,90)(1080,90)(1080,106){31}
//: {32}(1064,95)(938,95){33}
//: {34}(936,93)(936,90)(950,90)(950,109){35}
//: {36}(934,95)(810,95){37}
//: {38}(808,93)(808,90)(823,90)(823,104){39}
//: {40}(806,95)(752,95)(752,95)(679,95){41}
//: {42}(677,93)(677,90)(689,90)(689,117){43}
//: {44}(675,95)(565,95){45}
//: {46}(561,95)(346,95){47}
//: {48}(342,95)(162,95)(162,81)(147,81)(147,91){49}
//: {50}(344,97)(344,100)(357,100)(357,116){51}
//: {52}(563,97)(563,107)(563,107)(563,113){53}
//: {54}(1365,97)(1365,110){55}
//: {56}(1477,97)(1477,112){57}
//: {58}(1621,97)(1621,116){59}
//: {60}(1733,97)(1733,115){61}
//: {62}(1881,97)(1881,107)(1883,107)(1883,123){63}
//: {64}(2016,97)(2016,123){65}
//: {66}(2131,97)(2131,107)(2133,107)(2133,122){67}
//: {68}(2270,97)(2270,107)(2272,107)(2272,121){69}
//: {70}(2397,97)(2397,128){71}
//: {72}(2536,97)(2536,107)(2535,107)(2535,133){73}
output Cout;    //: /sn:0 {0}(99,332)(-62,332)(-62,266)(16,266){1}
output [17:0] Out;    //: /sn:0 {0}(1294,662)(1294,622)(1341,622)(1341,607)(#:1331,607){1}
wire w32;    //: /sn:0 {0}(1508,295)(1508,285)(1534,285)(1534,339)(1560,339){1}
wire w6;    //: /sn:0 {0}(801,294)(801,208)(809,208)(809,193){1}
wire w7;    //: /sn:0 {0}(1203,382)(1203,406)(1263,406)(1263,486){1}
wire [8:0] w45;    //: /sn:0 {0}(#:1325,612)(1314,612)(1314,569)(1358,569)(#:1358,493){1}
wire w60;    //: /sn:0 {0}(2258,210)(2258,288)(2244,288)(2244,303){1}
wire w46;    //: /sn:0 {0}(1378,487)(1378,468)(2270,468)(2270,391){1}
wire w61;    //: /sn:0 {0}(2540,392)(2540,482)(1398,482)(1398,487){1}
wire w56;    //: /sn:0 {0}(2119,211)(2119,286)(2117,286)(2117,301){1}
wire w16;    //: /sn:0 {0}(1026,332)(1021,332)(1021,275)(981,275)(981,294){1}
wire w14;    //: /sn:0 {0}(470,336)(406,336)(406,281)(372,281)(372,294){1}
wire w89;    //: /sn:0 {0}(2111,38)(2111,46)(2113,46)(2113,122){1}
wire w15;    //: /sn:0 {0}(1351,199)(1351,279)(1319,279)(1319,294){1}
wire w19;    //: /sn:0 {0}(862,294)(862,263)(889,263)(889,336)(891,336){1}
wire w4;    //: /sn:0 {0}(635,294)(635,224)(675,224)(675,206){1}
wire w38;    //: /sn:0 {0}(1037,38)(1037,91)(1060,91)(1060,106){1}
wire w51;    //: /sn:0 {0}(2049,300)(2049,290)(2073,290)(2073,343)(2088,343){1}
wire w0;    //: /sn:0 {0}(1418,337)(1405,337)(1405,284)(1380,284)(1380,294){1}
wire w3;    //: /sn:0 {0}(154,378)(154,479)(1193,479)(1193,486){1}
wire w66;    //: /sn:0 {0}(1615,385)(1615,435)(1328,435)(1328,487){1}
wire w64;    //: /sn:0 {0}(2383,217)(2383,290)(2373,290)(2373,305){1}
wire w37;    //: /sn:0 {0}(1650,297)(1650,287)(1679,287)(1679,341)(1693,341){1}
wire w63;    //: /sn:0 {0}(2434,305)(2434,295)(2462,295)(2462,346)(2485,346){1}
wire w34;    //: /sn:0 {0}(917,38)(917,67)(930,67)(930,109){1}
wire w43;    //: /sn:0 {0}(1783,299)(1783,290)(1816,290)(1816,341)(1831,341){1}
wire w21;    //: /sn:0 {0}(1081,378)(1081,431)(1253,431)(1253,486){1}
wire [8:0] w76;    //: /sn:0 {0}(#:1233,492)(1233,602)(#:1325,602){1}
wire w54;    //: /sn:0 {0}(2014,388)(2014,458)(1358,458)(1358,487){1}
wire w58;    //: /sn:0 {0}(1886,387)(1886,452)(1348,452)(1348,487){1}
wire w31;    //: /sn:0 {0}(661,382)(661,461)(1223,461)(1223,486){1}
wire w28;    //: /sn:0 {0}(1189,197)(1189,248)(1177,248)(1177,294){1}
wire w36;    //: /sn:0 {0}(1473,383)(1473,413)(1318,413)(1318,487){1}
wire w24;    //: /sn:0 {0}(1055,290)(1055,280)(1066,280)(1066,195){1}
wire w23;    //: /sn:0 {0}(668,38)(668,67)(669,67)(669,117){1}
wire w20;    //: /sn:0 {0}(544,38)(544,55)(543,55)(543,113){1}
wire w41;    //: /sn:0 {0}(1155,38)(1155,39)(1183,39)(1183,108){1}
wire w1;    //: /sn:0 {0}(128,290)(128,254)(133,254)(133,180){1}
wire w25;    //: /sn:0 {0}(1238,294)(1238,284)(1265,284)(1265,336)(1290,336){1}
wire w98;    //: /sn:0 {0}(2510,38)(2510,46)(2515,46)(2515,133){1}
wire w74;    //: /sn:0 {0}(1455,38)(1455,46)(1457,46)(1457,112){1}
wire w92;    //: /sn:0 {0}(2254,38)(2254,46)(2252,46)(2252,121){1}
wire w18;    //: /sn:0 {0}(920,294)(920,213)(936,213)(936,198){1}
wire w8;    //: /sn:0 {0}(772,336)(720,336)(720,261)(696,261)(696,294){1}
wire w35;    //: /sn:0 {0}(946,382)(946,437)(1243,437)(1243,486){1}
wire w71;    //: /sn:0 {0}(1345,110)(1345,38){1}
wire w68;    //: /sn:0 {0}(2521,222)(2521,289)(2514,289)(2514,304){1}
wire w30;    //: /sn:0 {0}(827,382)(827,454)(1233,454)(1233,486){1}
wire w22;    //: /sn:0 {0}(1148,336)(1147,336)(1147,261)(1116,261)(1116,290){1}
wire w17;    //: /sn:0 {0}(334,38)(334,70)(337,70)(337,116){1}
wire w59;    //: /sn:0 {0}(2305,303)(2305,287)(2334,287)(2334,345){1}
//: {2}(2336,347)(2344,347){3}
//: {4}(2332,347)(2327,347){5}
wire w62;    //: /sn:0 {0}(1748,387)(1748,446)(1338,446)(1338,487){1}
wire w44;    //: /sn:0 {0}(1719,204)(1719,284)(1722,284)(1722,299){1}
wire w2;    //: /sn:0 {0}(606,336)(584,336)(584,239)(560,239)(560,294){1}
wire w12;    //: /sn:0 {0}(105,38)(105,74)(127,74)(127,91){1}
wire w49;    //: /sn:0 {0}(525,382)(525,466)(1213,466)(1213,486){1}
wire w83;    //: /sn:0 {0}(1863,38)(1863,123){1}
wire w77;    //: /sn:0 {0}(1599,38)(1599,46)(1601,46)(1601,116){1}
wire w10;    //: /sn:0 {0}(1345,382)(1345,410)(1273,410)(1273,486){1}
wire w13;    //: /sn:0 {0}(282,336)(228,336)(228,268)(189,268)(189,290){1}
wire w27;    //: /sn:0 {0}(785,38)(785,94)(803,94)(803,104){1}
wire w95;    //: /sn:0 {0}(2370,38)(2370,46)(2377,46)(2377,128){1}
wire w86;    //: /sn:0 {0}(1996,38)(1996,123){1}
wire w52;    //: /sn:0 {0}(2002,212)(2002,285)(1988,285)(1988,300){1}
wire w48;    //: /sn:0 {0}(1869,212)(1869,284)(1860,284)(1860,299){1}
wire w33;    //: /sn:0 {0}(1463,201)(1463,280)(1447,280)(1447,295){1}
wire w5;    //: /sn:0 {0}(311,294)(311,289)(343,289)(343,205){1}
wire w80;    //: /sn:0 {0}(1715,38)(1715,46)(1713,46)(1713,115){1}
wire w47;    //: /sn:0 {0}(1921,299)(1921,286)(1949,286)(1949,340){1}
//: {2}(1951,342)(1959,342){3}
//: {4}(1947,342)(1942,342){5}
wire w29;    //: /sn:0 {0}(337,382)(337,473)(1203,473)(1203,486){1}
wire w50;    //: /sn:0 {0}(1368,487)(1368,463)(2143,463)(2143,389){1}
wire w42;    //: /sn:0 {0}(1388,487)(1388,473)(2399,473)(2399,393){1}
wire w9;    //: /sn:0 {0}(499,294)(499,289)(549,289)(549,202){1}
wire w55;    //: /sn:0 {0}(2178,301)(2178,276)(2212,276)(2212,345)(2215,345){1}
wire w39;    //: /sn:0 {0}(1607,205)(1607,271)(1589,271)(1589,297){1}
//: enddecls

  //: joint g61 (minus) @(1881, 95) /w:[ 15 -1 16 62 ]
  //: IN g4 (In) @(44,34) /sn:0 /w:[ 37 ]
  myEXOR g8 (.A(minus), .B(w17), .Out(w5));   //: @(313, 117) /sz:(60, 87) /R:3 /sn:0 /p:[ Ti0>51 Ti1>1 Bo0<1 ]
  //: joint g58 (minus) @(1477, 95) /w:[ 21 -1 22 56 ]
  myEXOR g55 (.A(minus), .B(w98), .Out(w68));   //: @(2491, 134) /sz:(60, 87) /R:3 /sn:0 /p:[ Ti0>73 Ti1>1 Bo0<0 ]
  myEXOR g51 (.A(minus), .B(w86), .Out(w52));   //: @(1972, 124) /sz:(60, 87) /R:3 /sn:0 /p:[ Ti0>65 Ti1>1 Bo0<0 ]
  MyHA g37 (.B(w33), .A(w32), .cout(w0), .S(w36));   //: @(1419, 296) /sz:(107, 86) /sn:0 /p:[ Ti0>1 Ti1>0 Lo0<0 Bo0<0 ]
  assign w12 = In[17]; //: TAP g13 @(105,32) /sn:0 /R:1 /w:[ 0 36 35 ] /ss:1
  MyHA g3 (.A(w8), .B(w4), .cout(w2), .S(w31));   //: @(607, 295) /sz:(107, 86) /sn:0 /p:[ Ti0>1 Ti1>0 Lo0<0 Bo0<0 ]
  assign w38 = In[11]; //: TAP g34 @(1037,32) /sn:0 /R:1 /w:[ 0 24 23 ] /ss:1
  assign w98 = In[0]; //: TAP g76 @(2510,32) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  //: joint g65 (minus) @(2397, 95) /w:[ 7 -1 8 70 ]
  MyHA g2 (.A(w2), .B(w9), .cout(w14), .S(w49));   //: @(471, 295) /sz:(107, 86) /sn:0 /p:[ Ti0>1 Ti1>0 Lo0<0 Bo0<0 ]
  assign w45 = {w36, w66, w62, w58, w54, w50, w46, w42, w61}; //: CONCAT g77  @(1358,492) /sn:0 /R:3 /w:[ 1 1 1 1 1 1 0 0 0 1 ] /dr:1 /tp:0 /drp:1
  //: joint g59 (minus) @(1621, 95) /w:[ 19 -1 20 58 ]
  assign w86 = In[4]; //: TAP g72 @(1996,32) /sn:0 /R:1 /w:[ 0 10 9 ] /ss:1
  MyHA g1 (.A(w14), .B(w5), .cout(w13), .S(w29));   //: @(283, 295) /sz:(107, 86) /sn:0 /p:[ Ti0>1 Ti1>0 Lo0<0 Bo0<0 ]
  //: joint g64 (minus) @(2270, 95) /w:[ 9 -1 10 68 ]
  //: joint g16 (minus) @(563, 95) /w:[ 45 -1 46 52 ]
  assign w23 = In[14]; //: TAP g11 @(668,32) /sn:0 /R:1 /w:[ 0 30 29 ] /ss:1
  myEXOR g50 (.A(minus), .B(w83), .Out(w48));   //: @(1839, 124) /sz:(60, 87) /R:3 /sn:0 /p:[ Ti0>63 Ti1>1 Bo0<0 ]
  myEXOR g10 (.A(minus), .B(w23), .Out(w4));   //: @(645, 118) /sz:(60, 87) /R:3 /sn:0 /p:[ Ti0>43 Ti1>1 Bo0<1 ]
  //: joint g28 (minus) @(936, 95) /w:[ 33 34 36 -1 ]
  assign Out = {w76, w45}; //: CONCAT g78  @(1330,607) /sn:0 /w:[ 1 1 0 ] /dr:0 /tp:0 /drp:1
  myEXOR g27 (.A(minus), .B(w41), .Out(w28));   //: @(1159, 109) /sz:(60, 87) /R:3 /sn:0 /p:[ Ti0>27 Ti1>1 Bo0<0 ]
  assign w27 = In[13]; //: TAP g32 @(785,32) /sn:0 /R:1 /w:[ 0 28 27 ] /ss:1
  assign w76 = {w3, w29, w49, w31, w30, w35, w21, w7, w10}; //: CONCAT g19  @(1233,491) /sn:0 /R:3 /w:[ 0 1 1 1 1 1 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  assign w77 = In[7]; //: TAP g69 @(1599,32) /sn:0 /R:1 /w:[ 0 16 15 ] /ss:1
  MyHA g38 (.B(w39), .A(w37), .cout(w32), .S(w66));   //: @(1561, 298) /sz:(107, 86) /sn:0 /p:[ Ti0>1 Ti1>0 Lo0<1 Bo0<0 ]
  //: OUT g6 (Out) @(1294,659) /sn:0 /R:3 /w:[ 0 ]
  assign w95 = In[1]; //: TAP g75 @(2370,32) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  //: joint g57 (minus) @(1365, 95) /w:[ 23 -1 24 54 ]
  myEXOR g53 (.A(minus), .B(w92), .Out(w60));   //: @(2228, 122) /sz:(60, 87) /R:3 /sn:0 /p:[ Ti0>69 Ti1>1 Bo0<0 ]
  myEXOR g9 (.A(minus), .B(w20), .Out(w9));   //: @(519, 114) /sz:(60, 87) /R:3 /sn:0 /p:[ Ti0>53 Ti1>1 Bo0<1 ]
  myEXOR g7 (.A(minus), .B(w12), .Out(w1));   //: @(103, 92) /sz:(60, 87) /R:3 /sn:0 /p:[ Ti0>49 Ti1>1 Bo0<1 ]
  assign w83 = In[5]; //: TAP g71 @(1863,32) /sn:0 /R:1 /w:[ 0 12 11 ] /ss:1
  //: joint g15 (w47) @(1949, 342) /w:[ 2 1 4 -1 ]
  //: joint g31 (minus) @(1188, 95) /w:[ 25 26 28 -1 ]
  MyHA g20 (.B(w6), .A(w19), .cout(w8), .S(w30));   //: @(773, 295) /sz:(107, 86) /sn:0 /p:[ Ti0>0 Ti1>0 Lo0<0 Bo0<0 ]
  assign w74 = In[8]; //: TAP g68 @(1455,32) /sn:0 /R:1 /w:[ 0 18 17 ] /ss:1
  assign w71 = In[9]; //: TAP g67 @(1345,32) /sn:0 /R:1 /w:[ 1 20 19 ] /ss:1
  MyHA g39 (.B(w44), .A(w43), .cout(w37), .S(w62));   //: @(1694, 300) /sz:(107, 86) /sn:0 /p:[ Ti0>1 Ti1>0 Lo0<1 Bo0<0 ]
  myEXOR g48 (.A(minus), .B(w77), .Out(w39));   //: @(1577, 117) /sz:(60, 87) /R:3 /sn:0 /p:[ Ti0>59 Ti1>1 Bo0<0 ]
  MyHA g43 (.B(w60), .A(w59), .cout(w55), .S(w46));   //: @(2216, 304) /sz:(107, 86) /sn:0 /p:[ Ti0>1 Ti1>0 Lo0<1 Bo0<1 ]
  assign w89 = In[3]; //: TAP g73 @(2111,32) /sn:0 /R:1 /w:[ 0 8 7 ] /ss:1
  //: joint g62 (minus) @(2016, 95) /w:[ 13 -1 14 64 ]
  //: joint g29 (minus) @(808, 95) /w:[ 37 38 40 -1 ]
  myEXOR g25 (.A(minus), .B(w34), .Out(w18));   //: @(906, 110) /sz:(60, 87) /R:3 /sn:0 /p:[ Ti0>35 Ti1>1 Bo0<1 ]
  //: joint g17 (minus) @(344, 95) /w:[ 47 -1 48 50 ]
  //: joint g63 (minus) @(2131, 95) /w:[ 11 -1 12 66 ]
  myEXOR g52 (.A(minus), .B(w89), .Out(w56));   //: @(2089, 123) /sz:(60, 87) /R:3 /sn:0 /p:[ Ti0>67 Ti1>1 Bo0<0 ]
  MyHA g42 (.B(w56), .A(w55), .cout(w51), .S(w50));   //: @(2089, 302) /sz:(107, 86) /sn:0 /p:[ Ti0>1 Ti1>0 Lo0<1 Bo0<1 ]
  assign w92 = In[2]; //: TAP g74 @(2254,32) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:1
  //: joint g56 (w59) @(2334, 347) /w:[ 2 1 4 -1 ]
  assign w20 = In[15]; //: TAP g14 @(544,32) /sn:0 /R:1 /w:[ 0 32 31 ] /ss:1
  //: IN g5 (minus) @(2591,28) /sn:0 /R:3 /w:[ 3 ]
  myEXOR g47 (.A(minus), .B(w74), .Out(w33));   //: @(1433, 113) /sz:(60, 87) /R:3 /sn:0 /p:[ Ti0>57 Ti1>1 Bo0<0 ]
  MyHA g44 (.B(w64), .A(w63), .cout(w59), .S(w42));   //: @(2345, 306) /sz:(107, 86) /sn:0 /p:[ Ti0>1 Ti1>0 Lo0<3 Bo0<1 ]
  //: joint g79 (minus) @(2576, 95) /w:[ 2 -1 4 1 ]
  //: OUT g80 (Cout) @(13,266) /sn:0 /w:[ 1 ]
  //: joint g36 (minus) @(677, 95) /w:[ 41 42 44 -1 ]
  myEXOR g24 (.A(minus), .B(w27), .Out(w6));   //: @(779, 105) /sz:(60, 87) /R:3 /sn:0 /p:[ Ti0>39 Ti1>1 Bo0<1 ]
  MyHA g21 (.B(w18), .A(w16), .cout(w19), .S(w35));   //: @(892, 295) /sz:(107, 86) /sn:0 /p:[ Ti0>0 Ti1>1 Lo0<1 Bo0<0 ]
  MyHA g41 (.B(w52), .A(w51), .cout(w47), .S(w54));   //: @(1960, 301) /sz:(107, 86) /sn:0 /p:[ Ti0>1 Ti1>0 Lo0<3 Bo0<0 ]
  MyHA g23 (.B(w28), .A(w25), .cout(w22), .S(w7));   //: @(1149, 295) /sz:(107, 86) /sn:0 /p:[ Ti0>1 Ti1>0 Lo0<0 Bo0<0 ]
  //: joint g60 (minus) @(1733, 95) /w:[ 17 -1 18 60 ]
  myEXOR g54 (.A(minus), .B(w95), .Out(w64));   //: @(2353, 129) /sz:(60, 87) /R:3 /sn:0 /p:[ Ti0>71 Ti1>1 Bo0<0 ]
  MyHA g40 (.B(w48), .A(w47), .cout(w43), .S(w58));   //: @(1832, 300) /sz:(107, 86) /sn:0 /p:[ Ti0>1 Ti1>0 Lo0<1 Bo0<0 ]
  assign w80 = In[6]; //: TAP g70 @(1715,32) /sn:0 /R:1 /w:[ 0 14 13 ] /ss:1
  myEXOR g46 (.A(minus), .B(w71), .Out(w15));   //: @(1321, 111) /sz:(60, 87) /R:3 /sn:0 /p:[ Ti0>55 Ti1>0 Bo0<0 ]
  MyHA g45 (.B(w68), .A(minus), .cout(w63), .S(w61));   //: @(2486, 305) /sz:(107, 86) /sn:0 /p:[ Ti0>1 Ti1>0 Lo0<1 Bo0<0 ]
  myEXOR g26 (.A(minus), .B(w38), .Out(w24));   //: @(1036, 107) /sz:(60, 87) /R:3 /sn:0 /p:[ Ti0>31 Ti1>1 Bo0<1 ]
  MyHA g22 (.B(w24), .A(w22), .cout(w16), .S(w21));   //: @(1027, 291) /sz:(107, 86) /sn:0 /p:[ Ti0>0 Ti1>1 Lo0<0 Bo0<0 ]
  MyHA g0 (.A(w13), .B(w1), .cout(Cout), .S(w3));   //: @(100, 291) /sz:(107, 86) /sn:0 /p:[ Ti0>1 Ti1>0 Lo0<0 Bo0<0 ]
  assign w41 = In[10]; //: TAP g35 @(1155,32) /sn:0 /R:1 /w:[ 0 22 21 ] /ss:1
  //: joint g66 (minus) @(2536, 95) /w:[ 5 -1 6 72 ]
  MyHA g18 (.B(w15), .A(w0), .cout(w25), .S(w10));   //: @(1291, 295) /sz:(107, 86) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<0 ]
  assign w17 = In[16]; //: TAP g12 @(334,32) /sn:0 /R:1 /w:[ 0 34 33 ] /ss:1
  //: joint g30 (minus) @(1066, 95) /w:[ 29 30 32 -1 ]
  assign w34 = In[12]; //: TAP g33 @(917,32) /sn:0 /R:1 /w:[ 0 26 25 ] /ss:1
  myEXOR g49 (.A(minus), .B(w80), .Out(w44));   //: @(1689, 116) /sz:(60, 87) /R:3 /sn:0 /p:[ Ti0>61 Ti1>1 Bo0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin myEXOR
module myEXOR(B, Out, A);
//: interface  /sz:(87, 60) /bd:[ Li0>B(36/60) Li1>A(16/60) Ro0<Out(30/60) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input B;    //: /sn:0 {0}(64,244)(122,244){1}
//: {2}(126,244)(395,244)(395,129)(408,129){3}
//: {4}(124,246)(124,353)(182,353){5}
input A;    //: /sn:0 {0}(51,95)(161,95){1}
//: {2}(165,95)(182,95)(182,67)(195,67){3}
//: {4}(163,97)(163,320)(422,320){5}
output Out;    //: /sn:0 {0}(690,198)(820,198){1}
wire w4;    //: /sn:0 {0}(422,348)(249,348)(249,371)(234,371){1}
wire w0;    //: /sn:0 {0}(247,85)(357,85)(357,101)(408,101){1}
wire w2;    //: /sn:0 {0}(500,116)(583,116)(583,183)(598,183){1}
wire w5;    //: /sn:0 {0}(514,335)(583,335)(583,211)(598,211){1}
//: enddecls

  myINV g4 (.In(B), .Out(w4));   //: @(183, 341) /sz:(50, 46) /sn:0 /p:[ Li0>5 Ro0<1 ]
  //: joint g8 (A) @(163, 95) /w:[ 2 -1 1 4 ]
  myINV g3 (.In(A), .Out(w0));   //: @(196, 55) /sz:(50, 46) /sn:0 /p:[ Li0>3 Ro0<0 ]
  myNAND2 g2 (.B(w5), .A(w2), .Out(Out));   //: @(599, 162) /sz:(90, 66) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]
  myNAND2 g1 (.B(w4), .A(A), .Out(w5));   //: @(423, 299) /sz:(90, 66) /sn:0 /p:[ Li0>0 Li1>5 Ro0<0 ]
  //: IN g6 (B) @(62,244) /sn:0 /w:[ 0 ]
  //: OUT g7 (Out) @(817,198) /sn:0 /w:[ 1 ]
  //: joint g9 (B) @(124, 244) /w:[ 2 -1 1 4 ]
  //: IN g5 (A) @(49,95) /sn:0 /w:[ 0 ]
  myNAND2 g0 (.B(B), .A(w0), .Out(w2));   //: @(409, 80) /sz:(90, 66) /sn:0 /p:[ Li0>3 Li1>1 Ro0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin MYREGISTER18
module MYREGISTER18(Clk, out, in);
//: interface  /sz:(123, 41) /bd:[ Li0>Clk(34/41) Li1>in[17:0](11/41) Ro0<out[17:0](12/41) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [17:0] in;    //: /sn:0 {0}(#:51,-6)(51,20){1}
//: {2}(51,21)(51,122){3}
//: {4}(51,123)(51,252){5}
//: {6}(51,253)(51,352){7}
//: {8}(51,353)(51,458){9}
//: {10}(51,459)(51,592){11}
//: {12}(51,593)(51,726){13}
//: {14}(51,727)(51,846){15}
//: {16}(51,847)(51,952){17}
//: {18}(51,953)(51,1052){19}
//: {20}(51,1053)(51,1161){21}
//: {22}(51,1162)(51,1287){23}
//: {24}(51,1288)(51,1400){25}
//: {26}(51,1401)(51,1514){27}
//: {28}(51,1515)(51,1613){29}
//: {30}(51,1614)(51,1723){31}
//: {32}(51,1724)(51,1826){33}
//: {34}(51,1827)(51,1964){35}
//: {36}(51,1965)(51,2083)(58,2083){37}
output [17:0] out;    //: /sn:0 {0}(#:938,818)(979,818)(979,817)(994,817){1}
input Clk;    //: /sn:0 {0}(450,2037)(450,2062)(385,2062)(385,2035)(139,2035){1}
//: {2}(137,2033)(137,1923){3}
//: {4}(139,1921)(446,1921)(446,1902){5}
//: {6}(137,1919)(137,1808){7}
//: {8}(139,1806)(450,1806)(450,1797){9}
//: {10}(137,1804)(137,1694){11}
//: {12}(139,1692)(456,1692)(456,1682){13}
//: {14}(137,1690)(137,1592){15}
//: {16}(139,1590)(463,1590)(463,1581){17}
//: {18}(137,1588)(137,1478){19}
//: {20}(139,1476)(464,1476)(464,1464){21}
//: {22}(137,1474)(137,1365){23}
//: {24}(139,1363)(465,1363)(465,1349){25}
//: {26}(137,1361)(137,1244){27}
//: {28}(139,1242)(468,1242)(468,1230){29}
//: {30}(137,1240)(137,1136){31}
//: {32}(139,1134)(473,1134)(473,1118){33}
//: {34}(137,1132)(137,1014){35}
//: {36}(139,1012)(391,1012)(391,1030)(476,1030)(476,1021){37}
//: {38}(137,1010)(137,926){39}
//: {40}(139,924)(480,924)(480,910){41}
//: {42}(137,922)(137,833){43}
//: {44}(139,831)(421,831)(421,812)(479,812)(479,794){45}
//: {46}(137,829)(137,698){47}
//: {48}(139,696)(479,696)(479,663){49}
//: {50}(137,694)(137,558){51}
//: {52}(139,556)(479,556)(479,535){53}
//: {54}(137,554)(137,439){55}
//: {56}(139,437)(479,437)(479,413){57}
//: {58}(137,435)(137,331){59}
//: {60}(139,329)(478,329)(478,308){61}
//: {62}(137,327)(137,228){63}
//: {64}(139,226)(391,226)(391,208)(478,208)(478,193){65}
//: {66}(137,224)(137,89)(478,89)(478,83){67}
//: {68}(137,2037)(137,2067)(132,2067){69}
wire w32;    //: /sn:0 {0}(506,1731)(612,1731)(612,1338)(745,1338){1}
wire w6;    //: /sn:0 {0}(429,243)(63,243)(63,253)(55,253){1}
wire w7;    //: /sn:0 {0}(532,955)(725,955)(725,511)(699,511)(699,496)(709,496){1}
wire w16;    //: /sn:0 {0}(529,1052)(730,1052)(730,1278)(745,1278){1}
wire w14;    //: /sn:0 {0}(535,469)(623,469)(623,456)(709,456){1}
wire w4;    //: /sn:0 {0}(407,1617)(63,1617)(63,1614)(55,1614){1}
wire w19;    //: /sn:0 {0}(419,1165)(63,1165)(63,1162)(55,1162){1}
wire w15;    //: /sn:0 {0}(430,598)(63,598)(63,593)(55,593){1}
wire w0;    //: /sn:0 {0}(429,18)(63,18)(63,21)(55,21){1}
wire w3;    //: /sn:0 {0}(429,128)(63,128)(63,123)(55,123){1}
wire w37;    //: /sn:0 {0}(401,1972)(63,1972)(63,1965)(55,1965){1}
wire w34;    //: /sn:0 {0}(397,1837)(63,1837)(63,1827)(55,1827){1}
wire w21;    //: /sn:0 {0}(431,845)(63,845)(63,847)(55,847){1}
wire w31;    //: /sn:0 {0}(414,1516)(63,1516)(63,1515)(55,1515){1}
wire w28;    //: /sn:0 {0}(415,1399)(63,1399)(63,1401)(55,1401){1}
wire w36;    //: /sn:0 {0}(502,1836)(628,1836)(628,1348)(745,1348){1}
wire w24;    //: /sn:0 {0}(524,1164)(670,1164)(670,1288)(745,1288){1}
wire w20;    //: /sn:0 {0}(535,728)(669,728)(669,476)(709,476){1}
wire w23;    //: /sn:0 {0}(709,486)(704,486)(704,844)(536,844){1}
wire w1;    //: /sn:0 {0}(427,956)(63,956)(63,953)(55,953){1}
wire w25;    //: /sn:0 {0}(416,1284)(63,1284)(63,1288)(55,1288){1}
wire [8:0] w35;    //: /sn:0 {0}(#:751,1318)(917,1318)(917,823)(932,823){1}
wire w8;    //: /sn:0 {0}(709,436)(616,436)(616,242)(534,242){1}
wire w18;    //: /sn:0 {0}(430,729)(63,729)(63,727)(55,727){1}
wire w30;    //: /sn:0 {0}(520,1398)(523,1398)(523,1308)(745,1308){1}
wire w22;    //: /sn:0 {0}(512,1616)(588,1616)(588,1328)(745,1328){1}
wire w17;    //: /sn:0 {0}(535,597)(656,597)(656,466)(709,466){1}
wire w2;    //: /sn:0 {0}(709,416)(702,416)(702,17)(534,17){1}
wire w11;    //: /sn:0 {0}(709,446)(550,446)(550,347)(535,347){1}
wire w12;    //: /sn:0 {0}(430,470)(63,470)(63,459)(55,459){1}
wire w10;    //: /sn:0 {0}(424,1053)(55,1053){1}
wire [8:0] w13;    //: /sn:0 {0}(#:715,456)(917,456)(917,813)(932,813){1}
wire w27;    //: /sn:0 {0}(521,1283)(551,1283)(551,1298)(745,1298){1}
wire w33;    //: /sn:0 {0}(745,1318)(534,1318)(534,1515)(519,1515){1}
wire w5;    //: /sn:0 {0}(709,426)(644,426)(644,127)(534,127){1}
wire w9;    //: /sn:0 {0}(430,348)(63,348)(63,353)(55,353){1}
wire w39;    //: /sn:0 {0}(506,1971)(672,1971)(672,1358)(745,1358){1}
wire w26;    //: /sn:0 {0}(401,1732)(63,1732)(63,1724)(55,1724){1}
//: enddecls

  FlipFlopDet g4 (.D(w12), .Clk(Clk), .Y(w14));   //: @(431, 449) /sz:(103, 85) /sn:0 /p:[ Li0>0 Bi0>53 Ro0<0 ]
  //: IN g8 (Clk) @(130,2067) /sn:0 /w:[ 69 ]
  //: OUT g58 (out) @(991,817) /sn:0 /w:[ 1 ]
  assign w37 = in[17]; //: TAP g55 @(49,1965) /sn:0 /R:2 /w:[ 1 36 35 ] /ss:1
  assign w34 = in[16]; //: TAP g51 @(49,1827) /sn:0 /R:2 /w:[ 1 34 33 ] /ss:1
  //: joint g37 (Clk) @(137, 1134) /w:[ 32 34 -1 31 ]
  assign w10 = in[9]; //: TAP g34 @(49,1053) /sn:0 /R:2 /w:[ 1 20 19 ] /ss:1
  FlipFlopDet g3 (.D(w9), .Clk(Clk), .Y(w11));   //: @(431, 327) /sz:(103, 85) /sn:0 /p:[ Li0>0 Bi0>57 Ro0<1 ]
  //: joint g13 (Clk) @(137, 696) /w:[ 48 50 -1 47 ]
  FlipFlopDet g2 (.D(w6), .Clk(Clk), .Y(w8));   //: @(430, 222) /sz:(103, 85) /sn:0 /p:[ Li0>0 Bi0>61 Ro0<1 ]
  FlipFlopDet g1 (.D(w3), .Clk(Clk), .Y(w5));   //: @(430, 107) /sz:(103, 85) /sn:0 /p:[ Li0>0 Bi0>65 Ro0<1 ]
  //: joint g11 (Clk) @(137, 437) /w:[ 56 58 -1 55 ]
  //: IN g16 (in) @(51,-8) /sn:0 /R:3 /w:[ 0 ]
  assign w26 = in[15]; //: TAP g50 @(49,1724) /sn:0 /R:2 /w:[ 1 32 31 ] /ss:1
  FlipFlopDet g28 (.D(w10), .Clk(Clk), .Y(w16));   //: @(425, 1032) /sz:(103, 85) /sn:0 /p:[ Li0>0 Bi0>33 Ro0<0 ]
  //: joint g10 (Clk) @(137, 329) /w:[ 60 62 -1 59 ]
  FlipFlopDet g32 (.D(w31), .Clk(Clk), .Y(w33));   //: @(415, 1495) /sz:(103, 85) /sn:0 /p:[ Li0>0 Bi0>17 Ro0<1 ]
  FlipFlopDet g27 (.D(w1), .Clk(Clk), .Y(w7));   //: @(428, 935) /sz:(103, 85) /sn:0 /p:[ Li0>0 Bi0>37 Ro0<0 ]
  assign w6 = in[2]; //: TAP g19 @(49,253) /sn:0 /R:2 /w:[ 1 6 5 ] /ss:1
  //: joint g38 (Clk) @(137, 1242) /w:[ 28 30 -1 27 ]
  FlipFlopDet g6 (.D(w18), .Clk(Clk), .Y(w20));   //: @(431, 708) /sz:(103, 85) /sn:0 /p:[ Li0>0 Bi0>45 Ro0<0 ]
  assign w35 = {w39, w36, w32, w22, w33, w30, w27, w24, w16}; //: CONCAT g57  @(750,1318) /sn:0 /w:[ 0 1 1 1 1 0 1 1 1 1 ] /dr:1 /tp:0 /drp:1
  //: joint g53 (Clk) @(137, 1806) /w:[ 8 10 -1 7 ]
  FlipFlopDet g7 (.D(w21), .Clk(Clk), .Y(w23));   //: @(432, 824) /sz:(103, 85) /sn:0 /p:[ Li0>0 Bi0>41 Ro0<1 ]
  //: joint g9 (Clk) @(137, 226) /w:[ 64 66 -1 63 ]
  FlipFlopDet g31 (.D(w28), .Clk(Clk), .Y(w30));   //: @(416, 1378) /sz:(103, 85) /sn:0 /p:[ Li0>0 Bi0>21 Ro0<0 ]
  //: joint g15 (Clk) @(137, 924) /w:[ 40 42 -1 39 ]
  assign w9 = in[3]; //: TAP g20 @(49,353) /sn:0 /R:2 /w:[ 1 8 7 ] /ss:1
  assign w25 = in[11]; //: TAP g39 @(49,1288) /sn:0 /R:2 /w:[ 1 24 23 ] /ss:1
  FlipFlopDet g48 (.D(w37), .Clk(Clk), .Y(w39));   //: @(402, 1951) /sz:(103, 85) /sn:0 /p:[ Li0>0 Bi0>0 Ro0<0 ]
  assign w31 = in[13]; //: TAP g43 @(49,1515) /sn:0 /R:2 /w:[ 1 28 27 ] /ss:1
  assign out = {w35, w13}; //: CONCAT g25  @(937,818) /sn:0 /w:[ 0 1 1 ] /dr:1 /tp:0 /drp:1
  FlipFlopDet g29 (.D(w19), .Clk(Clk), .Y(w24));   //: @(420, 1144) /sz:(103, 85) /sn:0 /p:[ Li0>0 Bi0>29 Ro0<0 ]
  assign w0 = in[0]; //: TAP g17 @(49,21) /sn:0 /R:2 /w:[ 1 2 1 ] /ss:1
  //: joint g52 (Clk) @(137, 1692) /w:[ 12 14 -1 11 ]
  //: joint g42 (Clk) @(137, 1476) /w:[ 20 22 -1 19 ]
  //: joint g56 (Clk) @(137, 2035) /w:[ 1 2 -1 68 ]
  FlipFlopDet g5 (.D(w15), .Clk(Clk), .Y(w17));   //: @(431, 577) /sz:(103, 85) /sn:0 /p:[ Li0>0 Bi0>49 Ro0<0 ]
  //: joint g14 (Clk) @(137, 831) /w:[ 44 46 -1 43 ]
  FlipFlopDet g47 (.D(w34), .Clk(Clk), .Y(w36));   //: @(398, 1816) /sz:(103, 85) /sn:0 /p:[ Li0>0 Bi0>5 Ro0<0 ]
  //: joint g44 (Clk) @(137, 1590) /w:[ 16 18 -1 15 ]
  //: joint g36 (Clk) @(137, 1012) /w:[ 36 38 -1 35 ]
  assign w12 = in[4]; //: TAP g21 @(49,459) /sn:0 /R:2 /w:[ 1 10 9 ] /ss:1
  assign w21 = in[7]; //: TAP g24 @(49,847) /sn:0 /R:2 /w:[ 1 16 15 ] /ss:1
  assign w28 = in[12]; //: TAP g41 @(49,1401) /sn:0 /R:2 /w:[ 1 26 25 ] /ss:1
  assign w18 = in[6]; //: TAP g23 @(49,727) /sn:0 /R:2 /w:[ 1 14 13 ] /ss:1
  //: joint g54 (Clk) @(137, 1921) /w:[ 4 6 -1 3 ]
  //: joint g40 (Clk) @(137, 1363) /w:[ 24 26 -1 23 ]
  FlipFlopDet g46 (.D(w26), .Clk(Clk), .Y(w32));   //: @(402, 1711) /sz:(103, 85) /sn:0 /p:[ Li0>0 Bi0>9 Ro0<0 ]
  FlipFlopDet g45 (.D(w4), .Clk(Clk), .Y(w22));   //: @(408, 1596) /sz:(103, 85) /sn:0 /p:[ Li0>0 Bi0>13 Ro0<0 ]
  assign w19 = in[10]; //: TAP g35 @(49,1162) /sn:0 /R:2 /w:[ 1 22 21 ] /ss:1
  FlipFlopDet g0 (.D(w0), .Clk(Clk), .Y(w2));   //: @(430, -3) /sz:(103, 85) /sn:0 /p:[ Li0>0 Bi0>67 Ro0<1 ]
  assign w15 = in[5]; //: TAP g22 @(49,593) /sn:0 /R:2 /w:[ 1 12 11 ] /ss:1
  assign w13 = {w7, w23, w20, w17, w14, w11, w8, w5, w2}; //: CONCAT g26  @(714,456) /sn:0 /w:[ 0 1 0 1 1 1 0 0 0 0 ] /dr:1 /tp:0 /drp:1
  //: joint g12 (Clk) @(137, 556) /w:[ 52 54 -1 51 ]
  assign w3 = in[1]; //: TAP g18 @(49,123) /sn:0 /R:2 /w:[ 1 4 3 ] /ss:1
  assign w1 = in[8]; //: TAP g33 @(49,953) /sn:0 /R:2 /w:[ 1 18 17 ] /ss:1
  FlipFlopDet g30 (.D(w25), .Clk(Clk), .Y(w27));   //: @(417, 1263) /sz:(103, 85) /sn:0 /p:[ Li0>0 Bi0>25 Ro0<0 ]
  assign w4 = in[14]; //: TAP g49 @(49,1614) /sn:0 /R:2 /w:[ 1 30 29 ] /ss:1

endmodule
//: /netlistEnd

//: /netlistBegin FlipFlopDet
module FlipFlopDet(Clk, Y, D);
//: interface  /sz:(103, 85) /bd:[ Li0>D(21/85) Bi0>Clk(48/103) Ro0<Y(20/85) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input Clk;    //: /sn:0 {0}(408,387)(477,387)(477,301){1}
//: {2}(477,297)(477,230){3}
//: {4}(475,299)(429,299)(429,305)(386,305){5}
input D;    //: /sn:0 {0}(91,149)(202,149)(202,159)(217,159){1}
output Y;    //: /sn:0 {0}(613,151)(547,151)(547,154)(532,154){1}
wire w1;    //: /sn:0 {0}(280,232)(280,287)(334,287){1}
wire w2;    //: /sn:0 {0}(335,156)(399,156)(399,157)(414,157){1}
//: enddecls

  //: IN g4 (Clk) @(406,387) /sn:0 /w:[ 0 ]
  //: OUT g3 (Y) @(610,151) /sn:0 /w:[ 0 ]
  //: IN g2 (D) @(89,149) /sn:0 /w:[ 0 ]
  FlipFlopDLS g1 (.D(w2), .Clk(Clk), .Y(Y));   //: @(415, 133) /sz:(116, 96) /sn:0 /p:[ Li0>1 Bi0>3 Ro0<1 ]
  //: joint g6 (Clk) @(477, 299) /w:[ -1 2 4 1 ]
  myINV g5 (.In(Clk), .Out(w1));   //: @(335, 271) /sz:(50, 46) /R:2 /sn:0 /p:[ Ri0>5 Lo0<1 ]
  FlipFlopDLS g0 (.D(D), .Clk(w1), .Y(w2));   //: @(218, 135) /sz:(116, 96) /sn:0 /p:[ Li0>1 Bi0>0 Ro0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin myNOR
module myNOR(out, in2, in1);
//: interface  /sz:(117, 91) /bd:[ Li0>in2(70/91) Li1>in1(29/91) Ro0<out(47/91) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output out;    //: /sn:0 {0}(373,187)(373,215){1}
//: {2}(375,217)(385,217)(385,218)(517,218){3}
//: {4}(373,219)(373,245){5}
//: {6}(375,247)(438,247)(438,262){7}
//: {8}(371,247)(330,247)(330,265){9}
input in1;    //: /sn:0 {0}(176,129)(242,129)(242,128)(341,128){1}
//: {2}(343,126)(343,120)(360,120){3}
//: {4}(343,130)(343,270)(424,270){5}
supply1 w12;    //: /sn:0 {0}(373,61)(373,97)(374,97)(374,112){1}
input in2;    //: /sn:0 {0}(173,222)(299,222){1}
//: {2}(301,220)(301,178)(359,178){3}
//: {4}(301,224)(301,273)(316,273){5}
supply0 w13;    //: /sn:0 {0}(394,321)(394,300)(392,300)(392,296){1}
//: {2}(394,294)(438,294)(438,279){3}
//: {4}(390,294)(330,294)(330,282){5}
wire w0;    //: /sn:0 {0}(374,129)(374,155)(373,155)(373,170){1}
//: enddecls

  //: OUT g8 (out) @(514,218) /sn:0 /w:[ 3 ]
  //: VDD g4 (w12) @(384,61) /sn:0 /w:[ 0 ]
  //: joint g13 (in2) @(301, 222) /w:[ -1 2 1 4 ]
  _GGNMOS #(2, 1) g3 (.Z(out), .S(w13), .G(in1));   //: @(432,270) /sn:0 /w:[ 7 3 5 ]
  _GGNMOS #(2, 1) g2 (.Z(out), .S(w13), .G(in2));   //: @(324,273) /sn:0 /w:[ 9 5 5 ]
  _GGPMOS #(2, 1) g1 (.Z(out), .S(w0), .G(in2));   //: @(367,178) /sn:0 /w:[ 0 1 3 ]
  //: IN g11 (in2) @(171,222) /sn:0 /w:[ 0 ]
  //: IN g10 (in1) @(174,129) /sn:0 /w:[ 0 ]
  //: joint g6 (out) @(373, 247) /w:[ 6 5 8 -1 ]
  //: joint g9 (out) @(373, 217) /w:[ 2 1 -1 4 ]
  //: joint g7 (w13) @(392, 294) /w:[ 2 -1 4 1 ]
  //: GROUND g5 (w13) @(394,327) /sn:0 /w:[ 0 ]
  _GGPMOS #(2, 1) g0 (.Z(w0), .S(w12), .G(in1));   //: @(368,120) /sn:0 /w:[ 0 1 3 ]
  //: joint g12 (in1) @(343, 128) /w:[ -1 2 1 4 ]

endmodule
//: /netlistEnd

//: /netlistBegin MYREGISTER8
module MYREGISTER8(Clk, in, out);
//: interface  /sz:(88, 106) /bd:[ Li0>in[7:0](29/106) Li1>Clk(90/106) Ro0<out[7:0](33/106) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [7:0] in;    //: /sn:0 {0}(#:51,-6)(51,20){1}
//: {2}(51,21)(51,122){3}
//: {4}(51,123)(51,252){5}
//: {6}(51,253)(51,352){7}
//: {8}(51,353)(51,458){9}
//: {10}(51,459)(51,592){11}
//: {12}(51,593)(51,726){13}
//: {14}(51,727)(51,846){15}
//: {16}(51,847)(51,1040)(43,1040){17}
output [7:0] out;    //: /sn:0 {0}(#:715,456)(808,456){1}
input Clk;    //: /sn:0 {0}(480,910)(480,924)(139,924){1}
//: {2}(137,922)(137,833){3}
//: {4}(139,831)(421,831)(421,812)(479,812)(479,794){5}
//: {6}(137,829)(137,698){7}
//: {8}(139,696)(479,696)(479,663){9}
//: {10}(137,694)(137,558){11}
//: {12}(139,556)(479,556)(479,535){13}
//: {14}(137,554)(137,439){15}
//: {16}(139,437)(479,437)(479,413){17}
//: {18}(137,435)(137,331){19}
//: {20}(139,329)(478,329)(478,308){21}
//: {22}(137,327)(137,228){23}
//: {24}(139,226)(391,226)(391,208)(478,208)(478,193){25}
//: {26}(137,224)(137,89)(478,89)(478,83){27}
//: {28}(137,926)(137,1016)(127,1016){29}
wire w6;    //: /sn:0 {0}(429,243)(63,243)(63,253)(55,253){1}
wire w14;    //: /sn:0 {0}(535,469)(623,469)(623,461)(709,461){1}
wire w15;    //: /sn:0 {0}(430,598)(63,598)(63,593)(55,593){1}
wire w0;    //: /sn:0 {0}(429,18)(63,18)(63,21)(55,21){1}
wire w3;    //: /sn:0 {0}(429,128)(63,128)(63,123)(55,123){1}
wire w21;    //: /sn:0 {0}(431,845)(63,845)(63,847)(55,847){1}
wire w20;    //: /sn:0 {0}(535,728)(669,728)(669,481)(709,481){1}
wire w23;    //: /sn:0 {0}(709,491)(704,491)(704,844)(536,844){1}
wire w8;    //: /sn:0 {0}(709,441)(616,441)(616,242)(534,242){1}
wire w18;    //: /sn:0 {0}(430,729)(63,729)(63,727)(55,727){1}
wire w17;    //: /sn:0 {0}(535,597)(656,597)(656,471)(709,471){1}
wire w2;    //: /sn:0 {0}(709,421)(702,421)(702,17)(534,17){1}
wire w11;    //: /sn:0 {0}(709,451)(550,451)(550,347)(535,347){1}
wire w12;    //: /sn:0 {0}(430,470)(63,470)(63,459)(55,459){1}
wire w5;    //: /sn:0 {0}(709,431)(644,431)(644,127)(534,127){1}
wire w9;    //: /sn:0 {0}(430,348)(63,348)(63,353)(55,353){1}
//: enddecls

  FlipFlopDet g4 (.D(w12), .Clk(Clk), .Y(w14));   //: @(431, 449) /sz:(103, 85) /sn:0 /p:[ Li0>0 Bi0>13 Ro0<0 ]
  //: IN g8 (Clk) @(125,1016) /sn:0 /w:[ 29 ]
  FlipFlopDet g3 (.D(w9), .Clk(Clk), .Y(w11));   //: @(431, 327) /sz:(103, 85) /sn:0 /p:[ Li0>0 Bi0>17 Ro0<1 ]
  //: joint g13 (Clk) @(137, 696) /w:[ 8 10 -1 7 ]
  FlipFlopDet g2 (.D(w6), .Clk(Clk), .Y(w8));   //: @(430, 222) /sz:(103, 85) /sn:0 /p:[ Li0>0 Bi0>21 Ro0<1 ]
  FlipFlopDet g1 (.D(w3), .Clk(Clk), .Y(w5));   //: @(430, 107) /sz:(103, 85) /sn:0 /p:[ Li0>0 Bi0>25 Ro0<1 ]
  //: joint g11 (Clk) @(137, 437) /w:[ 16 18 -1 15 ]
  //: IN g16 (in) @(51,-8) /sn:0 /R:3 /w:[ 0 ]
  //: joint g10 (Clk) @(137, 329) /w:[ 20 22 -1 19 ]
  assign w6 = in[2]; //: TAP g19 @(49,253) /sn:0 /R:2 /w:[ 1 6 5 ] /ss:1
  FlipFlopDet g6 (.D(w18), .Clk(Clk), .Y(w20));   //: @(431, 708) /sz:(103, 85) /sn:0 /p:[ Li0>0 Bi0>5 Ro0<0 ]
  FlipFlopDet g7 (.D(w21), .Clk(Clk), .Y(w23));   //: @(432, 824) /sz:(103, 85) /sn:0 /p:[ Li0>0 Bi0>0 Ro0<1 ]
  //: joint g9 (Clk) @(137, 226) /w:[ 24 26 -1 23 ]
  //: joint g15 (Clk) @(137, 924) /w:[ 1 2 -1 28 ]
  assign w9 = in[3]; //: TAP g20 @(49,353) /sn:0 /R:2 /w:[ 1 8 7 ] /ss:1
  assign w0 = in[0]; //: TAP g17 @(49,21) /sn:0 /R:2 /w:[ 1 2 1 ] /ss:1
  //: OUT g25 (out) @(805,456) /sn:0 /w:[ 1 ]
  FlipFlopDet g5 (.D(w15), .Clk(Clk), .Y(w17));   //: @(431, 577) /sz:(103, 85) /sn:0 /p:[ Li0>0 Bi0>9 Ro0<0 ]
  //: joint g14 (Clk) @(137, 831) /w:[ 4 6 -1 3 ]
  assign w12 = in[4]; //: TAP g21 @(49,459) /sn:0 /R:2 /w:[ 1 10 9 ] /ss:1
  assign w21 = in[7]; //: TAP g24 @(49,847) /sn:0 /R:2 /w:[ 1 16 15 ] /ss:1
  assign w18 = in[6]; //: TAP g23 @(49,727) /sn:0 /R:2 /w:[ 1 14 13 ] /ss:1
  FlipFlopDet g0 (.D(w0), .Clk(Clk), .Y(w2));   //: @(430, -3) /sz:(103, 85) /sn:0 /p:[ Li0>0 Bi0>27 Ro0<1 ]
  assign w15 = in[5]; //: TAP g22 @(49,593) /sn:0 /R:2 /w:[ 1 12 11 ] /ss:1
  assign out = {w23, w20, w17, w14, w11, w8, w5, w2}; //: CONCAT g26  @(714,456) /sn:0 /w:[ 0 0 1 1 1 0 0 0 0 ] /dr:1 /tp:0 /drp:1
  //: joint g12 (Clk) @(137, 556) /w:[ 12 14 -1 11 ]
  assign w3 = in[1]; //: TAP g18 @(49,123) /sn:0 /R:2 /w:[ 1 4 3 ] /ss:1

endmodule
//: /netlistEnd

//: /netlistBegin myINV
module myINV(Out, In);
//: interface  /sz:(50, 46) /bd:[ Li0>In(12/46) Ro0<Out(30/46) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input In;    //: /sn:0 {0}(369,203)(456,203){1}
//: {2}(458,201)(458,167)(487,167){3}
//: {4}(458,205)(458,250)(487,250){5}
supply1 w0;    //: /sn:0 {0}(501,159)(501,83){1}
supply0 w1;    //: /sn:0 {0}(501,341)(501,259){1}
output Out;    //: /sn:0 {0}(501,242)(501,204){1}
//: {2}(503,202)(618,202)(618,201)(621,201){3}
//: {4}(501,200)(501,176){5}
//: enddecls

  _GGPMOS #(2, 1) g4 (.Z(Out), .S(w0), .G(In));   //: @(495,167) /sn:0 /w:[ 5 0 3 ]
  //: GROUND g3 (w1) @(501,347) /sn:0 /w:[ 0 ]
  //: VDD g2 (w0) @(512,83) /sn:0 /w:[ 1 ]
  //: OUT g1 (Out) @(618,201) /sn:0 /w:[ 3 ]
  //: joint g6 (In) @(458, 203) /w:[ -1 2 1 4 ]
  //: joint g7 (Out) @(501, 202) /w:[ 2 4 -1 1 ]
  _GGNMOS #(2, 1) g5 (.Z(Out), .S(w1), .G(In));   //: @(495,250) /sn:0 /w:[ 0 1 5 ]
  //: IN g0 (In) @(367,203) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin FA
module FA(Cout, B, S, Cin, A);
//: interface  /sz:(90, 88) /bd:[ Ti0>A(22/90) Ti1>B(66/90) Ri0>Cin(38/88) Lo0<Cout(37/88) Bo0<S(46/90) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input B;    //: /sn:0 {0}(109,311)(234,311)(234,163)(249,163){1}
input A;    //: /sn:0 {0}(102,123)(234,123)(234,102)(249,102){1}
output Cout;    //: /sn:0 {0}(813,258)(878,258)(878,254)(938,254){1}
input Cin;    //: /sn:0 {0}(116,347)(428,347)(428,332)(443,332){1}
output S;    //: /sn:0 {0}(531,306)(832,306){1}
wire w4;    //: /sn:0 {0}(684,186)(746,186)(746,240)(761,240){1}
wire w3;    //: /sn:0 {0}(337,137)(428,137)(428,271)(443,271){1}
wire w0;    //: /sn:0 {0}(291,192)(291,202)(448,202)(448,168)(565,168){1}
wire w1;    //: /sn:0 {0}(485,361)(485,374)(552,374)(552,209)(565,209){1}
//: enddecls

  //: OUT g8 (Cout) @(935,254) /sn:0 /w:[ 1 ]
  myINV g3 (.In(w4), .Out(Cout));   //: @(762, 228) /sz:(50, 46) /sn:0 /p:[ Li0>1 Ro0<0 ]
  myNOR g2 (.in2(w1), .in1(w0), .out(w4));   //: @(566, 139) /sz:(117, 91) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]
  MyHA g1 (.A(w3), .B(Cin), .cout(w1), .S(S));   //: @(444, 254) /sz:(86, 107) /R:1 /sn:0 /p:[ Li0>1 Li1>1 Bo0<0 Ro0<0 ]
  //: IN g6 (B) @(107,311) /sn:0 /w:[ 0 ]
  //: OUT g9 (S) @(829,306) /sn:0 /w:[ 1 ]
  //: IN g7 (Cin) @(114,347) /sn:0 /w:[ 0 ]
  //: IN g5 (A) @(100,123) /sn:0 /w:[ 0 ]
  MyHA g0 (.A(A), .B(B), .cout(w0), .S(w3));   //: @(250, 85) /sz:(86, 107) /R:1 /sn:0 /p:[ Li0>1 Li1>1 Bo0<0 Ro0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin myNAND2
module myNAND2(Out, A, B);
//: interface  /sz:(90, 66) /bd:[ Li0>B(49/66) Li1>A(21/66) Ro0<Out(36/66) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input B;    //: /sn:0 {0}(210,323)(478,323){1}
//: {2}(482,323)(508,323){3}
//: {4}(480,321)(480,141)(544,141){5}
input A;    //: /sn:0 {0}(231,188)(409,188){1}
//: {2}(413,188)(431,188)(431,143)(444,143){3}
//: {4}(411,190)(411,249)(508,249){5}
output Out;    //: /sn:0 {0}(522,241)(522,211){1}
//: {2}(524,209)(749,209){3}
//: {4}(522,207)(522,167){5}
//: {6}(524,165)(558,165)(558,150){7}
//: {8}(520,165)(458,165)(458,152){9}
supply1 w12;    //: /sn:0 {0}(510,51)(510,116){1}
//: {2}(512,118)(558,118)(558,133){3}
//: {4}(508,118)(458,118)(458,135){5}
supply0 w13;    //: /sn:0 {0}(522,404)(522,332){1}
wire w6;    //: /sn:0 {0}(522,315)(522,258){1}
//: enddecls

  //: VDD g4 (w12) @(521,51) /sn:0 /w:[ 0 ]
  //: OUT g8 (Out) @(746,209) /sn:0 /w:[ 3 ]
  _GGNMOS #(2, 1) g3 (.Z(Out), .S(w6), .G(A));   //: @(516,249) /sn:0 /w:[ 0 1 5 ]
  //: joint g13 (B) @(480, 323) /w:[ 2 4 1 -1 ]
  _GGNMOS #(2, 1) g2 (.Z(w6), .S(w13), .G(B));   //: @(516,323) /sn:0 /w:[ 0 1 3 ]
  _GGPMOS #(2, 1) g1 (.Z(Out), .S(w12), .G(B));   //: @(552,141) /sn:0 /w:[ 7 3 5 ]
  //: joint g11 (Out) @(522, 209) /w:[ 2 4 -1 1 ]
  //: joint g10 (w12) @(510, 118) /w:[ 2 1 4 -1 ]
  //: IN g6 (A) @(229,188) /sn:0 /w:[ 0 ]
  //: IN g7 (B) @(208,323) /sn:0 /w:[ 0 ]
  //: joint g9 (Out) @(522, 165) /w:[ 6 -1 8 5 ]
  //: GROUND g5 (w13) @(522,410) /sn:0 /w:[ 0 ]
  _GGPMOS #(2, 1) g0 (.Z(Out), .S(w12), .G(A));   //: @(452,143) /sn:0 /w:[ 9 5 3 ]
  //: joint g12 (A) @(411, 188) /w:[ 2 -1 1 4 ]

endmodule
//: /netlistEnd

